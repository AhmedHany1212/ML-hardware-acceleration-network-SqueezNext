module BIAS_layer9_19_7 #(parameter N_adder_tree=16)(q);
output wire [N_adder_tree*18-1:0] q;


BIAS #(.value(18'b000000000100011000))  U0 (.q(q[18*(0+1)-1:18*0]));
BIAS #(.value(18'b000011001000011000))  U1 (.q(q[18*(1+1)-1:18*1]));
BIAS #(.value(18'b000000101010100100))  U2 (.q(q[18*(2+1)-1:18*2]));
BIAS #(.value(18'b110111011100001000))  U3 (.q(q[18*(3+1)-1:18*3]));
BIAS #(.value(18'b000011011001010000))  U4 (.q(q[18*(4+1)-1:18*4]));
BIAS #(.value(18'b000001010110001100))  U5 (.q(q[18*(5+1)-1:18*5]));
BIAS #(.value(18'b000001110010001000))  U6 (.q(q[18*(6+1)-1:18*6]));
BIAS #(.value(18'b000010101000110000))  U7 (.q(q[18*(7+1)-1:18*7]));
BIAS #(.value(18'b111101011101110100))  U8 (.q(q[18*(8+1)-1:18*8]));
BIAS #(.value(18'b111101011110100100))  U9 (.q(q[18*(9+1)-1:18*9]));
BIAS #(.value(18'b000010010111000100))  U10 (.q(q[18*(10+1)-1:18*10]));
BIAS #(.value(18'b000010100111001100))  U11 (.q(q[18*(11+1)-1:18*11]));
BIAS #(.value(18'b000000101101101100))  U12 (.q(q[18*(12+1)-1:18*12]));
BIAS #(.value(18'b000110110001001100))  U13 (.q(q[18*(13+1)-1:18*13]));
BIAS #(.value(18'b000001011000010000))  U14 (.q(q[18*(14+1)-1:18*14]));
BIAS #(.value(18'b000000011100101100))  U15 (.q(q[18*(15+1)-1:18*15]));


endmodule
