module adder_2in_FP(
 input 	signed  [17:0] a,b,
 output signed 	[17:0] out
 );
 
assign out=a+b;
endmodule


