module CONV15 #(parameter N=256,parameter ADDR_WIDTH=1)(addr,clk,q);
input wire [ADDR_WIDTH-1:0] addr;
output wire [N*16-1:0] q ;
input clk;
W_ROM #(.FILENAME("conv15/CONV15_1.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U0 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv15/CONV15_2.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U1 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv15/CONV15_3.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U2 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv15/CONV15_4.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U3 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv15/CONV15_5.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U4 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv15/CONV15_6.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U5 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv15/CONV15_7.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U6 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv15/CONV15_8.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U7 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv15/CONV15_9.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U8 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv15/CONV15_10.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U9 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv15/CONV15_11.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U10 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv15/CONV15_12.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U11 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv15/CONV15_13.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U12 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv15/CONV15_14.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U13 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv15/CONV15_15.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U14 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv15/CONV15_16.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U15 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv15/CONV15_17.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U16 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv15/CONV15_18.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U17 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv15/CONV15_19.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U18 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv15/CONV15_20.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U19 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv15/CONV15_21.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U20 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv15/CONV15_22.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U21 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv15/CONV15_23.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U22 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv15/CONV15_24.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U23 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv15/CONV15_25.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U24 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv15/CONV15_26.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U25 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv15/CONV15_27.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U26 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv15/CONV15_28.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U27 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv15/CONV15_29.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U28 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv15/CONV15_30.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U29 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv15/CONV15_31.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U30 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv15/CONV15_32.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U31 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv15/CONV15_33.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U32 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv15/CONV15_34.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U33 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv15/CONV15_35.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U34 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv15/CONV15_36.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U35 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv15/CONV15_37.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U36 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv15/CONV15_38.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U37 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv15/CONV15_39.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U38 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv15/CONV15_40.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U39 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv15/CONV15_41.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U40 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv15/CONV15_42.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U41 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv15/CONV15_43.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U42 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv15/CONV15_44.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U43 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv15/CONV15_45.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U44 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv15/CONV15_46.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U45 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv15/CONV15_47.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U46 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv15/CONV15_48.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U47 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv15/CONV15_49.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U48 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv15/CONV15_50.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U49 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv15/CONV15_51.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U50 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv15/CONV15_52.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U51 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv15/CONV15_53.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U52 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv15/CONV15_54.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U53 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv15/CONV15_55.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U54 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv15/CONV15_56.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U55 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv15/CONV15_57.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U56 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv15/CONV15_58.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U57 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv15/CONV15_59.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U58 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv15/CONV15_60.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U59 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv15/CONV15_61.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U60 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv15/CONV15_62.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U61 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv15/CONV15_63.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U62 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv15/CONV15_64.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U63 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(63+1)-1:16*63])); 
W_ROM #(.FILENAME("conv15/CONV15_65.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U64 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(64+1)-1:16*64])); 
W_ROM #(.FILENAME("conv15/CONV15_66.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U65 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(65+1)-1:16*65])); 
W_ROM #(.FILENAME("conv15/CONV15_67.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U66 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(66+1)-1:16*66])); 
W_ROM #(.FILENAME("conv15/CONV15_68.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U67 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(67+1)-1:16*67])); 
W_ROM #(.FILENAME("conv15/CONV15_69.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U68 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(68+1)-1:16*68])); 
W_ROM #(.FILENAME("conv15/CONV15_70.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U69 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(69+1)-1:16*69])); 
W_ROM #(.FILENAME("conv15/CONV15_71.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U70 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(70+1)-1:16*70])); 
W_ROM #(.FILENAME("conv15/CONV15_72.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U71 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(71+1)-1:16*71])); 
W_ROM #(.FILENAME("conv15/CONV15_73.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U72 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(72+1)-1:16*72])); 
W_ROM #(.FILENAME("conv15/CONV15_74.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U73 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(73+1)-1:16*73])); 
W_ROM #(.FILENAME("conv15/CONV15_75.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U74 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(74+1)-1:16*74])); 
W_ROM #(.FILENAME("conv15/CONV15_76.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U75 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(75+1)-1:16*75])); 
W_ROM #(.FILENAME("conv15/CONV15_77.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U76 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(76+1)-1:16*76])); 
W_ROM #(.FILENAME("conv15/CONV15_78.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U77 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(77+1)-1:16*77])); 
W_ROM #(.FILENAME("conv15/CONV15_79.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U78 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(78+1)-1:16*78])); 
W_ROM #(.FILENAME("conv15/CONV15_80.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U79 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(79+1)-1:16*79])); 
W_ROM #(.FILENAME("conv15/CONV15_81.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U80 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(80+1)-1:16*80])); 
W_ROM #(.FILENAME("conv15/CONV15_82.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U81 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(81+1)-1:16*81])); 
W_ROM #(.FILENAME("conv15/CONV15_83.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U82 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(82+1)-1:16*82])); 
W_ROM #(.FILENAME("conv15/CONV15_84.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U83 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(83+1)-1:16*83])); 
W_ROM #(.FILENAME("conv15/CONV15_85.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U84 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(84+1)-1:16*84])); 
W_ROM #(.FILENAME("conv15/CONV15_86.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U85 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(85+1)-1:16*85])); 
W_ROM #(.FILENAME("conv15/CONV15_87.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U86 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(86+1)-1:16*86])); 
W_ROM #(.FILENAME("conv15/CONV15_88.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U87 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(87+1)-1:16*87])); 
W_ROM #(.FILENAME("conv15/CONV15_89.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U88 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(88+1)-1:16*88])); 
W_ROM #(.FILENAME("conv15/CONV15_90.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U89 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(89+1)-1:16*89])); 
W_ROM #(.FILENAME("conv15/CONV15_91.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U90 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(90+1)-1:16*90])); 
W_ROM #(.FILENAME("conv15/CONV15_92.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U91 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(91+1)-1:16*91])); 
W_ROM #(.FILENAME("conv15/CONV15_93.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U92 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(92+1)-1:16*92])); 
W_ROM #(.FILENAME("conv15/CONV15_94.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U93 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(93+1)-1:16*93])); 
W_ROM #(.FILENAME("conv15/CONV15_95.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U94 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(94+1)-1:16*94])); 
W_ROM #(.FILENAME("conv15/CONV15_96.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U95 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(95+1)-1:16*95])); 
W_ROM #(.FILENAME("conv15/CONV15_97.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U96 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(96+1)-1:16*96])); 
W_ROM #(.FILENAME("conv15/CONV15_98.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U97 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(97+1)-1:16*97])); 
W_ROM #(.FILENAME("conv15/CONV15_99.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U98 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(98+1)-1:16*98])); 
W_ROM #(.FILENAME("conv15/CONV15_100.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U99 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(99+1)-1:16*99])); 
W_ROM #(.FILENAME("conv15/CONV15_101.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U100 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(100+1)-1:16*100])); 
W_ROM #(.FILENAME("conv15/CONV15_102.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U101 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(101+1)-1:16*101])); 
W_ROM #(.FILENAME("conv15/CONV15_103.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U102 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(102+1)-1:16*102])); 
W_ROM #(.FILENAME("conv15/CONV15_104.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U103 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(103+1)-1:16*103])); 
W_ROM #(.FILENAME("conv15/CONV15_105.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U104 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(104+1)-1:16*104])); 
W_ROM #(.FILENAME("conv15/CONV15_106.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U105 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(105+1)-1:16*105])); 
W_ROM #(.FILENAME("conv15/CONV15_107.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U106 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(106+1)-1:16*106])); 
W_ROM #(.FILENAME("conv15/CONV15_108.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U107 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(107+1)-1:16*107])); 
W_ROM #(.FILENAME("conv15/CONV15_109.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U108 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(108+1)-1:16*108])); 
W_ROM #(.FILENAME("conv15/CONV15_110.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U109 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(109+1)-1:16*109])); 
W_ROM #(.FILENAME("conv15/CONV15_111.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U110 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(110+1)-1:16*110])); 
W_ROM #(.FILENAME("conv15/CONV15_112.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U111 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(111+1)-1:16*111])); 
W_ROM #(.FILENAME("conv15/CONV15_113.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U112 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(112+1)-1:16*112])); 
W_ROM #(.FILENAME("conv15/CONV15_114.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U113 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(113+1)-1:16*113])); 
W_ROM #(.FILENAME("conv15/CONV15_115.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U114 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(114+1)-1:16*114])); 
W_ROM #(.FILENAME("conv15/CONV15_116.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U115 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(115+1)-1:16*115])); 
W_ROM #(.FILENAME("conv15/CONV15_117.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U116 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(116+1)-1:16*116])); 
W_ROM #(.FILENAME("conv15/CONV15_118.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U117 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(117+1)-1:16*117])); 
W_ROM #(.FILENAME("conv15/CONV15_119.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U118 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(118+1)-1:16*118])); 
W_ROM #(.FILENAME("conv15/CONV15_120.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U119 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(119+1)-1:16*119])); 
W_ROM #(.FILENAME("conv15/CONV15_121.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U120 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(120+1)-1:16*120])); 
W_ROM #(.FILENAME("conv15/CONV15_122.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U121 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(121+1)-1:16*121])); 
W_ROM #(.FILENAME("conv15/CONV15_123.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U122 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(122+1)-1:16*122])); 
W_ROM #(.FILENAME("conv15/CONV15_124.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U123 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(123+1)-1:16*123])); 
W_ROM #(.FILENAME("conv15/CONV15_125.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U124 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(124+1)-1:16*124])); 
W_ROM #(.FILENAME("conv15/CONV15_126.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U125 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(125+1)-1:16*125])); 
W_ROM #(.FILENAME("conv15/CONV15_127.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U126 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(126+1)-1:16*126])); 
W_ROM #(.FILENAME("conv15/CONV15_128.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U127 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(127+1)-1:16*127])); 
W_ROM #(.FILENAME("conv15/CONV15_129.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U128 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(128+1)-1:16*128])); 
W_ROM #(.FILENAME("conv15/CONV15_130.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U129 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(129+1)-1:16*129])); 
W_ROM #(.FILENAME("conv15/CONV15_131.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U130 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(130+1)-1:16*130])); 
W_ROM #(.FILENAME("conv15/CONV15_132.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U131 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(131+1)-1:16*131])); 
W_ROM #(.FILENAME("conv15/CONV15_133.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U132 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(132+1)-1:16*132])); 
W_ROM #(.FILENAME("conv15/CONV15_134.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U133 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(133+1)-1:16*133])); 
W_ROM #(.FILENAME("conv15/CONV15_135.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U134 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(134+1)-1:16*134])); 
W_ROM #(.FILENAME("conv15/CONV15_136.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U135 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(135+1)-1:16*135])); 
W_ROM #(.FILENAME("conv15/CONV15_137.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U136 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(136+1)-1:16*136])); 
W_ROM #(.FILENAME("conv15/CONV15_138.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U137 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(137+1)-1:16*137])); 
W_ROM #(.FILENAME("conv15/CONV15_139.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U138 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(138+1)-1:16*138])); 
W_ROM #(.FILENAME("conv15/CONV15_140.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U139 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(139+1)-1:16*139])); 
W_ROM #(.FILENAME("conv15/CONV15_141.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U140 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(140+1)-1:16*140])); 
W_ROM #(.FILENAME("conv15/CONV15_142.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U141 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(141+1)-1:16*141])); 
W_ROM #(.FILENAME("conv15/CONV15_143.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U142 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(142+1)-1:16*142])); 
W_ROM #(.FILENAME("conv15/CONV15_144.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U143 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(143+1)-1:16*143])); 
W_ROM #(.FILENAME("conv15/CONV15_145.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U144 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(144+1)-1:16*144])); 
W_ROM #(.FILENAME("conv15/CONV15_146.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U145 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(145+1)-1:16*145])); 
W_ROM #(.FILENAME("conv15/CONV15_147.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U146 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(146+1)-1:16*146])); 
W_ROM #(.FILENAME("conv15/CONV15_148.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U147 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(147+1)-1:16*147])); 
W_ROM #(.FILENAME("conv15/CONV15_149.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U148 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(148+1)-1:16*148])); 
W_ROM #(.FILENAME("conv15/CONV15_150.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U149 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(149+1)-1:16*149])); 
W_ROM #(.FILENAME("conv15/CONV15_151.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U150 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(150+1)-1:16*150])); 
W_ROM #(.FILENAME("conv15/CONV15_152.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U151 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(151+1)-1:16*151])); 
W_ROM #(.FILENAME("conv15/CONV15_153.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U152 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(152+1)-1:16*152])); 
W_ROM #(.FILENAME("conv15/CONV15_154.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U153 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(153+1)-1:16*153])); 
W_ROM #(.FILENAME("conv15/CONV15_155.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U154 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(154+1)-1:16*154])); 
W_ROM #(.FILENAME("conv15/CONV15_156.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U155 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(155+1)-1:16*155])); 
W_ROM #(.FILENAME("conv15/CONV15_157.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U156 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(156+1)-1:16*156])); 
W_ROM #(.FILENAME("conv15/CONV15_158.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U157 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(157+1)-1:16*157])); 
W_ROM #(.FILENAME("conv15/CONV15_159.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U158 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(158+1)-1:16*158])); 
W_ROM #(.FILENAME("conv15/CONV15_160.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U159 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(159+1)-1:16*159])); 
W_ROM #(.FILENAME("conv15/CONV15_161.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U160 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(160+1)-1:16*160])); 
W_ROM #(.FILENAME("conv15/CONV15_162.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U161 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(161+1)-1:16*161])); 
W_ROM #(.FILENAME("conv15/CONV15_163.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U162 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(162+1)-1:16*162])); 
W_ROM #(.FILENAME("conv15/CONV15_164.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U163 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(163+1)-1:16*163])); 
W_ROM #(.FILENAME("conv15/CONV15_165.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U164 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(164+1)-1:16*164])); 
W_ROM #(.FILENAME("conv15/CONV15_166.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U165 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(165+1)-1:16*165])); 
W_ROM #(.FILENAME("conv15/CONV15_167.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U166 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(166+1)-1:16*166])); 
W_ROM #(.FILENAME("conv15/CONV15_168.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U167 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(167+1)-1:16*167])); 
W_ROM #(.FILENAME("conv15/CONV15_169.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U168 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(168+1)-1:16*168])); 
W_ROM #(.FILENAME("conv15/CONV15_170.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U169 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(169+1)-1:16*169])); 
W_ROM #(.FILENAME("conv15/CONV15_171.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U170 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(170+1)-1:16*170])); 
W_ROM #(.FILENAME("conv15/CONV15_172.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U171 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(171+1)-1:16*171])); 
W_ROM #(.FILENAME("conv15/CONV15_173.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U172 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(172+1)-1:16*172])); 
W_ROM #(.FILENAME("conv15/CONV15_174.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U173 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(173+1)-1:16*173])); 
W_ROM #(.FILENAME("conv15/CONV15_175.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U174 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(174+1)-1:16*174])); 
W_ROM #(.FILENAME("conv15/CONV15_176.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U175 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(175+1)-1:16*175])); 
W_ROM #(.FILENAME("conv15/CONV15_177.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U176 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(176+1)-1:16*176])); 
W_ROM #(.FILENAME("conv15/CONV15_178.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U177 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(177+1)-1:16*177])); 
W_ROM #(.FILENAME("conv15/CONV15_179.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U178 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(178+1)-1:16*178])); 
W_ROM #(.FILENAME("conv15/CONV15_180.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U179 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(179+1)-1:16*179])); 
W_ROM #(.FILENAME("conv15/CONV15_181.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U180 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(180+1)-1:16*180])); 
W_ROM #(.FILENAME("conv15/CONV15_182.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U181 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(181+1)-1:16*181])); 
W_ROM #(.FILENAME("conv15/CONV15_183.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U182 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(182+1)-1:16*182])); 
W_ROM #(.FILENAME("conv15/CONV15_184.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U183 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(183+1)-1:16*183])); 
W_ROM #(.FILENAME("conv15/CONV15_185.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U184 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(184+1)-1:16*184])); 
W_ROM #(.FILENAME("conv15/CONV15_186.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U185 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(185+1)-1:16*185])); 
W_ROM #(.FILENAME("conv15/CONV15_187.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U186 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(186+1)-1:16*186])); 
W_ROM #(.FILENAME("conv15/CONV15_188.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U187 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(187+1)-1:16*187])); 
W_ROM #(.FILENAME("conv15/CONV15_189.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U188 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(188+1)-1:16*188])); 
W_ROM #(.FILENAME("conv15/CONV15_190.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U189 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(189+1)-1:16*189])); 
W_ROM #(.FILENAME("conv15/CONV15_191.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U190 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(190+1)-1:16*190])); 
W_ROM #(.FILENAME("conv15/CONV15_192.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U191 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(191+1)-1:16*191])); 
W_ROM #(.FILENAME("conv15/CONV15_193.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U192 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(192+1)-1:16*192])); 
W_ROM #(.FILENAME("conv15/CONV15_194.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U193 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(193+1)-1:16*193])); 
W_ROM #(.FILENAME("conv15/CONV15_195.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U194 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(194+1)-1:16*194])); 
W_ROM #(.FILENAME("conv15/CONV15_196.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U195 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(195+1)-1:16*195])); 
W_ROM #(.FILENAME("conv15/CONV15_197.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U196 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(196+1)-1:16*196])); 
W_ROM #(.FILENAME("conv15/CONV15_198.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U197 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(197+1)-1:16*197])); 
W_ROM #(.FILENAME("conv15/CONV15_199.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U198 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(198+1)-1:16*198])); 
W_ROM #(.FILENAME("conv15/CONV15_200.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U199 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(199+1)-1:16*199])); 
W_ROM #(.FILENAME("conv15/CONV15_201.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U200 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(200+1)-1:16*200])); 
W_ROM #(.FILENAME("conv15/CONV15_202.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U201 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(201+1)-1:16*201])); 
W_ROM #(.FILENAME("conv15/CONV15_203.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U202 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(202+1)-1:16*202])); 
W_ROM #(.FILENAME("conv15/CONV15_204.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U203 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(203+1)-1:16*203])); 
W_ROM #(.FILENAME("conv15/CONV15_205.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U204 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(204+1)-1:16*204])); 
W_ROM #(.FILENAME("conv15/CONV15_206.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U205 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(205+1)-1:16*205])); 
W_ROM #(.FILENAME("conv15/CONV15_207.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U206 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(206+1)-1:16*206])); 
W_ROM #(.FILENAME("conv15/CONV15_208.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U207 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(207+1)-1:16*207])); 
W_ROM #(.FILENAME("conv15/CONV15_209.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U208 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(208+1)-1:16*208])); 
W_ROM #(.FILENAME("conv15/CONV15_210.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U209 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(209+1)-1:16*209])); 
W_ROM #(.FILENAME("conv15/CONV15_211.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U210 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(210+1)-1:16*210])); 
W_ROM #(.FILENAME("conv15/CONV15_212.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U211 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(211+1)-1:16*211])); 
W_ROM #(.FILENAME("conv15/CONV15_213.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U212 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(212+1)-1:16*212])); 
W_ROM #(.FILENAME("conv15/CONV15_214.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U213 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(213+1)-1:16*213])); 
W_ROM #(.FILENAME("conv15/CONV15_215.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U214 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(214+1)-1:16*214])); 
W_ROM #(.FILENAME("conv15/CONV15_216.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U215 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(215+1)-1:16*215])); 
W_ROM #(.FILENAME("conv15/CONV15_217.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U216 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(216+1)-1:16*216])); 
W_ROM #(.FILENAME("conv15/CONV15_218.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U217 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(217+1)-1:16*217])); 
W_ROM #(.FILENAME("conv15/CONV15_219.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U218 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(218+1)-1:16*218])); 
W_ROM #(.FILENAME("conv15/CONV15_220.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U219 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(219+1)-1:16*219])); 
W_ROM #(.FILENAME("conv15/CONV15_221.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U220 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(220+1)-1:16*220])); 
W_ROM #(.FILENAME("conv15/CONV15_222.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U221 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(221+1)-1:16*221])); 
W_ROM #(.FILENAME("conv15/CONV15_223.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U222 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(222+1)-1:16*222])); 
W_ROM #(.FILENAME("conv15/CONV15_224.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U223 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(223+1)-1:16*223])); 
W_ROM #(.FILENAME("conv15/CONV15_225.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U224 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(224+1)-1:16*224])); 
W_ROM #(.FILENAME("conv15/CONV15_226.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U225 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(225+1)-1:16*225])); 
W_ROM #(.FILENAME("conv15/CONV15_227.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U226 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(226+1)-1:16*226])); 
W_ROM #(.FILENAME("conv15/CONV15_228.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U227 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(227+1)-1:16*227])); 
W_ROM #(.FILENAME("conv15/CONV15_229.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U228 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(228+1)-1:16*228])); 
W_ROM #(.FILENAME("conv15/CONV15_230.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U229 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(229+1)-1:16*229])); 
W_ROM #(.FILENAME("conv15/CONV15_231.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U230 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(230+1)-1:16*230])); 
W_ROM #(.FILENAME("conv15/CONV15_232.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U231 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(231+1)-1:16*231])); 
W_ROM #(.FILENAME("conv15/CONV15_233.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U232 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(232+1)-1:16*232])); 
W_ROM #(.FILENAME("conv15/CONV15_234.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U233 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(233+1)-1:16*233])); 
W_ROM #(.FILENAME("conv15/CONV15_235.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U234 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(234+1)-1:16*234])); 
W_ROM #(.FILENAME("conv15/CONV15_236.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U235 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(235+1)-1:16*235])); 
W_ROM #(.FILENAME("conv15/CONV15_237.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U236 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(236+1)-1:16*236])); 
W_ROM #(.FILENAME("conv15/CONV15_238.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U237 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(237+1)-1:16*237])); 
W_ROM #(.FILENAME("conv15/CONV15_239.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U238 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(238+1)-1:16*238])); 
W_ROM #(.FILENAME("conv15/CONV15_240.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U239 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(239+1)-1:16*239])); 
W_ROM #(.FILENAME("conv15/CONV15_241.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U240 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(240+1)-1:16*240])); 
W_ROM #(.FILENAME("conv15/CONV15_242.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U241 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(241+1)-1:16*241])); 
W_ROM #(.FILENAME("conv15/CONV15_243.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U242 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(242+1)-1:16*242])); 
W_ROM #(.FILENAME("conv15/CONV15_244.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U243 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(243+1)-1:16*243])); 
W_ROM #(.FILENAME("conv15/CONV15_245.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U244 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(244+1)-1:16*244])); 
W_ROM #(.FILENAME("conv15/CONV15_246.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U245 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(245+1)-1:16*245])); 
W_ROM #(.FILENAME("conv15/CONV15_247.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U246 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(246+1)-1:16*246])); 
W_ROM #(.FILENAME("conv15/CONV15_248.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U247 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(247+1)-1:16*247])); 
W_ROM #(.FILENAME("conv15/CONV15_249.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U248 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(248+1)-1:16*248])); 
W_ROM #(.FILENAME("conv15/CONV15_250.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U249 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(249+1)-1:16*249])); 
W_ROM #(.FILENAME("conv15/CONV15_251.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U250 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(250+1)-1:16*250])); 
W_ROM #(.FILENAME("conv15/CONV15_252.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U251 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(251+1)-1:16*251])); 
W_ROM #(.FILENAME("conv15/CONV15_253.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U252 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(252+1)-1:16*252])); 
W_ROM #(.FILENAME("conv15/CONV15_254.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U253 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(253+1)-1:16*253])); 
W_ROM #(.FILENAME("conv15/CONV15_255.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U254 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(254+1)-1:16*254])); 
W_ROM #(.FILENAME("conv15/CONV15_256.txt"),.weight_addr_WIDTH(1),.NO_ROWS(2)) U255 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(255+1)-1:16*255])); 


endmodule
