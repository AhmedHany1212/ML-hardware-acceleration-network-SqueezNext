module BIAS_layer16_55_2 #(parameter N_adder_tree=16)(q);
output wire [N_adder_tree*18-1:0] q;


BIAS #(.value(18'b111010000100111100))  U0 (.q(q[18*(0+1)-1:18*0]));
BIAS #(.value(18'b111010110100010100))  U1 (.q(q[18*(1+1)-1:18*1]));
BIAS #(.value(18'b111011110100011000))  U2 (.q(q[18*(2+1)-1:18*2]));
BIAS #(.value(18'b000100001010010000))  U3 (.q(q[18*(3+1)-1:18*3]));
BIAS #(.value(18'b111010111001101100))  U4 (.q(q[18*(4+1)-1:18*4]));
BIAS #(.value(18'b111000101001101000))  U5 (.q(q[18*(5+1)-1:18*5]));
BIAS #(.value(18'b000011111001011000))  U6 (.q(q[18*(6+1)-1:18*6]));
BIAS #(.value(18'b000000110000011100))  U7 (.q(q[18*(7+1)-1:18*7]));
BIAS #(.value(18'b000000011000101100))  U8 (.q(q[18*(8+1)-1:18*8]));
BIAS #(.value(18'b111111110011011000))  U9 (.q(q[18*(9+1)-1:18*9]));
BIAS #(.value(18'b000100001100110100))  U10 (.q(q[18*(10+1)-1:18*10]));
BIAS #(.value(18'b000101010000111100))  U11 (.q(q[18*(11+1)-1:18*11]));
BIAS #(.value(18'b111101101110101000))  U12 (.q(q[18*(12+1)-1:18*12]));
BIAS #(.value(18'b111110100000010000))  U13 (.q(q[18*(13+1)-1:18*13]));
BIAS #(.value(18'b111001001010010000))  U14 (.q(q[18*(14+1)-1:18*14]));
BIAS #(.value(18'b001000010010001000))  U15 (.q(q[18*(15+1)-1:18*15]));


endmodule
