//we have 192 distributed rom each one has different 11 num(9 and 2 padding) so we need 192 num at time (192*16 bits)

module CONV1 #(parameter N_weight_out=192,parameter weight_addr_WIDTH=4)(weight_addr,clk,weight_out);
input wire [weight_addr_WIDTH-1:0] weight_addr;
input clk;
output wire [N_weight_out*16-1:0] weight_out ;
W_ROM #(.FILENAME("conv1/CONV1_1.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U0 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv1/CONV1_2.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U1 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv1/CONV1_3.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U2 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv1/CONV1_4.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U3 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv1/CONV1_5.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U4 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv1/CONV1_6.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U5 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv1/CONV1_7.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U6 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv1/CONV1_8.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U7 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv1/CONV1_9.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U8 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv1/CONV1_10.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U9 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv1/CONV1_11.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U10 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv1/CONV1_12.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U11 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv1/CONV1_13.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U12 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv1/CONV1_14.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U13 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv1/CONV1_15.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U14 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv1/CONV1_16.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U15 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv1/CONV1_17.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U16 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv1/CONV1_18.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U17 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv1/CONV1_19.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U18 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv1/CONV1_20.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U19 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv1/CONV1_21.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U20 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv1/CONV1_22.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U21 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv1/CONV1_23.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U22 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv1/CONV1_24.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U23 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv1/CONV1_25.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U24 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv1/CONV1_26.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U25 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv1/CONV1_27.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U26 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv1/CONV1_28.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U27 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv1/CONV1_29.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U28 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv1/CONV1_30.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U29 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv1/CONV1_31.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U30 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv1/CONV1_32.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U31 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv1/CONV1_33.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U32 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv1/CONV1_34.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U33 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv1/CONV1_35.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U34 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv1/CONV1_36.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U35 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv1/CONV1_37.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U36 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv1/CONV1_38.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U37 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv1/CONV1_39.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U38 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv1/CONV1_40.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U39 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv1/CONV1_41.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U40 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv1/CONV1_42.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U41 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv1/CONV1_43.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U42 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv1/CONV1_44.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U43 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv1/CONV1_45.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U44 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv1/CONV1_46.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U45 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv1/CONV1_47.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U46 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv1/CONV1_48.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U47 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv1/CONV1_49.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U48 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv1/CONV1_50.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U49 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv1/CONV1_51.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U50 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv1/CONV1_52.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U51 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv1/CONV1_53.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U52 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv1/CONV1_54.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U53 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv1/CONV1_55.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U54 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv1/CONV1_56.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U55 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv1/CONV1_57.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U56 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv1/CONV1_58.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U57 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv1/CONV1_59.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U58 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv1/CONV1_60.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U59 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv1/CONV1_61.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U60 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv1/CONV1_62.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U61 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv1/CONV1_63.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U62 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv1/CONV1_64.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U63 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(63+1)-1:16*63])); 
W_ROM #(.FILENAME("conv1/CONV1_65.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U64 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(64+1)-1:16*64])); 
W_ROM #(.FILENAME("conv1/CONV1_66.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U65 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(65+1)-1:16*65])); 
W_ROM #(.FILENAME("conv1/CONV1_67.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U66 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(66+1)-1:16*66])); 
W_ROM #(.FILENAME("conv1/CONV1_68.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U67 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(67+1)-1:16*67])); 
W_ROM #(.FILENAME("conv1/CONV1_69.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U68 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(68+1)-1:16*68])); 
W_ROM #(.FILENAME("conv1/CONV1_70.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U69 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(69+1)-1:16*69])); 
W_ROM #(.FILENAME("conv1/CONV1_71.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U70 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(70+1)-1:16*70])); 
W_ROM #(.FILENAME("conv1/CONV1_72.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U71 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(71+1)-1:16*71])); 
W_ROM #(.FILENAME("conv1/CONV1_73.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U72 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(72+1)-1:16*72])); 
W_ROM #(.FILENAME("conv1/CONV1_74.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U73 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(73+1)-1:16*73])); 
W_ROM #(.FILENAME("conv1/CONV1_75.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U74 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(74+1)-1:16*74])); 
W_ROM #(.FILENAME("conv1/CONV1_76.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U75 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(75+1)-1:16*75])); 
W_ROM #(.FILENAME("conv1/CONV1_77.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U76 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(76+1)-1:16*76])); 
W_ROM #(.FILENAME("conv1/CONV1_78.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U77 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(77+1)-1:16*77])); 
W_ROM #(.FILENAME("conv1/CONV1_79.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U78 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(78+1)-1:16*78])); 
W_ROM #(.FILENAME("conv1/CONV1_80.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U79 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(79+1)-1:16*79])); 
W_ROM #(.FILENAME("conv1/CONV1_81.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U80 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(80+1)-1:16*80])); 
W_ROM #(.FILENAME("conv1/CONV1_82.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U81 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(81+1)-1:16*81])); 
W_ROM #(.FILENAME("conv1/CONV1_83.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U82 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(82+1)-1:16*82])); 
W_ROM #(.FILENAME("conv1/CONV1_84.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U83 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(83+1)-1:16*83])); 
W_ROM #(.FILENAME("conv1/CONV1_85.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U84 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(84+1)-1:16*84])); 
W_ROM #(.FILENAME("conv1/CONV1_86.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U85 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(85+1)-1:16*85])); 
W_ROM #(.FILENAME("conv1/CONV1_87.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U86 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(86+1)-1:16*86])); 
W_ROM #(.FILENAME("conv1/CONV1_88.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U87 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(87+1)-1:16*87])); 
W_ROM #(.FILENAME("conv1/CONV1_89.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U88 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(88+1)-1:16*88])); 
W_ROM #(.FILENAME("conv1/CONV1_90.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U89 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(89+1)-1:16*89])); 
W_ROM #(.FILENAME("conv1/CONV1_91.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U90 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(90+1)-1:16*90])); 
W_ROM #(.FILENAME("conv1/CONV1_92.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U91 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(91+1)-1:16*91])); 
W_ROM #(.FILENAME("conv1/CONV1_93.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U92 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(92+1)-1:16*92])); 
W_ROM #(.FILENAME("conv1/CONV1_94.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U93 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(93+1)-1:16*93])); 
W_ROM #(.FILENAME("conv1/CONV1_95.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U94 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(94+1)-1:16*94])); 
W_ROM #(.FILENAME("conv1/CONV1_96.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U95 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(95+1)-1:16*95])); 
W_ROM #(.FILENAME("conv1/CONV1_97.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U96 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(96+1)-1:16*96])); 
W_ROM #(.FILENAME("conv1/CONV1_98.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U97 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(97+1)-1:16*97])); 
W_ROM #(.FILENAME("conv1/CONV1_99.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U98 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(98+1)-1:16*98])); 
W_ROM #(.FILENAME("conv1/CONV1_100.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U99 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(99+1)-1:16*99])); 
W_ROM #(.FILENAME("conv1/CONV1_101.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U100 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(100+1)-1:16*100])); 
W_ROM #(.FILENAME("conv1/CONV1_102.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U101 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(101+1)-1:16*101])); 
W_ROM #(.FILENAME("conv1/CONV1_103.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U102 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(102+1)-1:16*102])); 
W_ROM #(.FILENAME("conv1/CONV1_104.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U103 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(103+1)-1:16*103])); 
W_ROM #(.FILENAME("conv1/CONV1_105.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U104 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(104+1)-1:16*104])); 
W_ROM #(.FILENAME("conv1/CONV1_106.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U105 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(105+1)-1:16*105])); 
W_ROM #(.FILENAME("conv1/CONV1_107.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U106 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(106+1)-1:16*106])); 
W_ROM #(.FILENAME("conv1/CONV1_108.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U107 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(107+1)-1:16*107])); 
W_ROM #(.FILENAME("conv1/CONV1_109.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U108 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(108+1)-1:16*108])); 
W_ROM #(.FILENAME("conv1/CONV1_110.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U109 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(109+1)-1:16*109])); 
W_ROM #(.FILENAME("conv1/CONV1_111.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U110 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(110+1)-1:16*110])); 
W_ROM #(.FILENAME("conv1/CONV1_112.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U111 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(111+1)-1:16*111])); 
W_ROM #(.FILENAME("conv1/CONV1_113.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U112 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(112+1)-1:16*112])); 
W_ROM #(.FILENAME("conv1/CONV1_114.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U113 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(113+1)-1:16*113])); 
W_ROM #(.FILENAME("conv1/CONV1_115.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U114 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(114+1)-1:16*114])); 
W_ROM #(.FILENAME("conv1/CONV1_116.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U115 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(115+1)-1:16*115])); 
W_ROM #(.FILENAME("conv1/CONV1_117.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U116 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(116+1)-1:16*116])); 
W_ROM #(.FILENAME("conv1/CONV1_118.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U117 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(117+1)-1:16*117])); 
W_ROM #(.FILENAME("conv1/CONV1_119.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U118 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(118+1)-1:16*118])); 
W_ROM #(.FILENAME("conv1/CONV1_120.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U119 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(119+1)-1:16*119])); 
W_ROM #(.FILENAME("conv1/CONV1_121.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U120 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(120+1)-1:16*120])); 
W_ROM #(.FILENAME("conv1/CONV1_122.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U121 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(121+1)-1:16*121])); 
W_ROM #(.FILENAME("conv1/CONV1_123.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U122 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(122+1)-1:16*122])); 
W_ROM #(.FILENAME("conv1/CONV1_124.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U123 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(123+1)-1:16*123])); 
W_ROM #(.FILENAME("conv1/CONV1_125.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U124 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(124+1)-1:16*124])); 
W_ROM #(.FILENAME("conv1/CONV1_126.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U125 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(125+1)-1:16*125])); 
W_ROM #(.FILENAME("conv1/CONV1_127.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U126 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(126+1)-1:16*126])); 
W_ROM #(.FILENAME("conv1/CONV1_128.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U127 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(127+1)-1:16*127])); 
W_ROM #(.FILENAME("conv1/CONV1_129.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U128 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(128+1)-1:16*128])); 
W_ROM #(.FILENAME("conv1/CONV1_130.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U129 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(129+1)-1:16*129])); 
W_ROM #(.FILENAME("conv1/CONV1_131.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U130 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(130+1)-1:16*130])); 
W_ROM #(.FILENAME("conv1/CONV1_132.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U131 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(131+1)-1:16*131])); 
W_ROM #(.FILENAME("conv1/CONV1_133.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U132 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(132+1)-1:16*132])); 
W_ROM #(.FILENAME("conv1/CONV1_134.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U133 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(133+1)-1:16*133])); 
W_ROM #(.FILENAME("conv1/CONV1_135.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U134 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(134+1)-1:16*134])); 
W_ROM #(.FILENAME("conv1/CONV1_136.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U135 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(135+1)-1:16*135])); 
W_ROM #(.FILENAME("conv1/CONV1_137.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U136 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(136+1)-1:16*136])); 
W_ROM #(.FILENAME("conv1/CONV1_138.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U137 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(137+1)-1:16*137])); 
W_ROM #(.FILENAME("conv1/CONV1_139.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U138 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(138+1)-1:16*138])); 
W_ROM #(.FILENAME("conv1/CONV1_140.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U139 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(139+1)-1:16*139])); 
W_ROM #(.FILENAME("conv1/CONV1_141.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U140 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(140+1)-1:16*140])); 
W_ROM #(.FILENAME("conv1/CONV1_142.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U141 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(141+1)-1:16*141])); 
W_ROM #(.FILENAME("conv1/CONV1_143.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U142 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(142+1)-1:16*142])); 
W_ROM #(.FILENAME("conv1/CONV1_144.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U143 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(143+1)-1:16*143])); 
W_ROM #(.FILENAME("conv1/CONV1_145.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U144 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(144+1)-1:16*144])); 
W_ROM #(.FILENAME("conv1/CONV1_146.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U145 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(145+1)-1:16*145])); 
W_ROM #(.FILENAME("conv1/CONV1_147.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U146 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(146+1)-1:16*146])); 
W_ROM #(.FILENAME("conv1/CONV1_148.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U147 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(147+1)-1:16*147])); 
W_ROM #(.FILENAME("conv1/CONV1_149.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U148 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(148+1)-1:16*148])); 
W_ROM #(.FILENAME("conv1/CONV1_150.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U149 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(149+1)-1:16*149])); 
W_ROM #(.FILENAME("conv1/CONV1_151.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U150 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(150+1)-1:16*150])); 
W_ROM #(.FILENAME("conv1/CONV1_152.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U151 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(151+1)-1:16*151])); 
W_ROM #(.FILENAME("conv1/CONV1_153.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U152 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(152+1)-1:16*152])); 
W_ROM #(.FILENAME("conv1/CONV1_154.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U153 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(153+1)-1:16*153])); 
W_ROM #(.FILENAME("conv1/CONV1_155.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U154 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(154+1)-1:16*154])); 
W_ROM #(.FILENAME("conv1/CONV1_156.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U155 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(155+1)-1:16*155])); 
W_ROM #(.FILENAME("conv1/CONV1_157.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U156 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(156+1)-1:16*156])); 
W_ROM #(.FILENAME("conv1/CONV1_158.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U157 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(157+1)-1:16*157])); 
W_ROM #(.FILENAME("conv1/CONV1_159.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U158 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(158+1)-1:16*158])); 
W_ROM #(.FILENAME("conv1/CONV1_160.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U159 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(159+1)-1:16*159])); 
W_ROM #(.FILENAME("conv1/CONV1_161.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U160 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(160+1)-1:16*160])); 
W_ROM #(.FILENAME("conv1/CONV1_162.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U161 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(161+1)-1:16*161])); 
W_ROM #(.FILENAME("conv1/CONV1_163.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U162 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(162+1)-1:16*162])); 
W_ROM #(.FILENAME("conv1/CONV1_164.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U163 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(163+1)-1:16*163])); 
W_ROM #(.FILENAME("conv1/CONV1_165.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U164 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(164+1)-1:16*164])); 
W_ROM #(.FILENAME("conv1/CONV1_166.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U165 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(165+1)-1:16*165])); 
W_ROM #(.FILENAME("conv1/CONV1_167.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U166 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(166+1)-1:16*166])); 
W_ROM #(.FILENAME("conv1/CONV1_168.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U167 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(167+1)-1:16*167])); 
W_ROM #(.FILENAME("conv1/CONV1_169.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U168 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(168+1)-1:16*168])); 
W_ROM #(.FILENAME("conv1/CONV1_170.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U169 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(169+1)-1:16*169])); 
W_ROM #(.FILENAME("conv1/CONV1_171.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U170 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(170+1)-1:16*170])); 
W_ROM #(.FILENAME("conv1/CONV1_172.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U171 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(171+1)-1:16*171])); 
W_ROM #(.FILENAME("conv1/CONV1_173.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U172 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(172+1)-1:16*172])); 
W_ROM #(.FILENAME("conv1/CONV1_174.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U173 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(173+1)-1:16*173])); 
W_ROM #(.FILENAME("conv1/CONV1_175.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U174 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(174+1)-1:16*174])); 
W_ROM #(.FILENAME("conv1/CONV1_176.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U175 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(175+1)-1:16*175])); 
W_ROM #(.FILENAME("conv1/CONV1_177.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U176 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(176+1)-1:16*176])); 
W_ROM #(.FILENAME("conv1/CONV1_178.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U177 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(177+1)-1:16*177])); 
W_ROM #(.FILENAME("conv1/CONV1_179.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U178 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(178+1)-1:16*178])); 
W_ROM #(.FILENAME("conv1/CONV1_180.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U179 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(179+1)-1:16*179])); 
W_ROM #(.FILENAME("conv1/CONV1_181.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U180 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(180+1)-1:16*180])); 
W_ROM #(.FILENAME("conv1/CONV1_182.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U181 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(181+1)-1:16*181])); 
W_ROM #(.FILENAME("conv1/CONV1_183.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U182 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(182+1)-1:16*182])); 
W_ROM #(.FILENAME("conv1/CONV1_184.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U183 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(183+1)-1:16*183])); 
W_ROM #(.FILENAME("conv1/CONV1_185.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U184 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(184+1)-1:16*184])); 
W_ROM #(.FILENAME("conv1/CONV1_186.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U185 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(185+1)-1:16*185])); 
W_ROM #(.FILENAME("conv1/CONV1_187.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U186 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(186+1)-1:16*186])); 
W_ROM #(.FILENAME("conv1/CONV1_188.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U187 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(187+1)-1:16*187])); 
W_ROM #(.FILENAME("conv1/CONV1_189.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U188 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(188+1)-1:16*188])); 
W_ROM #(.FILENAME("conv1/CONV1_190.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U189 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(189+1)-1:16*189])); 
W_ROM #(.FILENAME("conv1/CONV1_191.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U190 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(190+1)-1:16*190])); 
W_ROM #(.FILENAME("conv1/CONV1_192.txt"),.weight_addr_WIDTH(4) ,.NO_ROWS(11)) U191 (.weight_addr(weight_addr), .clk(clk),.weight_out(weight_out[16*(191+1)-1:16*191])); 

endmodule
