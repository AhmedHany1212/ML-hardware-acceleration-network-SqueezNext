module BIAS_layer4 #(parameter N_adder_tree=8)(out,Z);
wire [16*18-1:0] q;
input wire Z;
output wire [N_adder_tree*18-1:0] out;
assign out= Z ? q[18*(7+1)-1:18*0] : q[18*(15+1)-1:18*8];

BIAS #(.value(18'b111111010000111000)) U0 (.q(q[18*(0+1)-1:18*0]));
BIAS #(.value(18'b111111111111010000)) U1 (.q(q[18*(1+1)-1:18*1])); 
BIAS #(.value(18'b000000000011110100)) U2 (.q(q[18*(2+1)-1:18*2]));
BIAS #(.value(18'b111111110010101100)) U3 (.q(q[18*(3+1)-1:18*3]));
BIAS #(.value(18'b111111011000111100)) U4 (.q(q[18*(4+1)-1:18*4])); 
BIAS #(.value(18'b000001000100001100)) U5 (.q(q[18*(5+1)-1:18*5])); 
BIAS #(.value(18'b000000001100110100)) U6 (.q(q[18*(6+1)-1:18*6])); 
BIAS #(.value(18'b000001101011000100)) U7 (.q(q[18*(7+1)-1:18*7])); 

BIAS #(.value(18'b000010001000111100)) U8  (.q(q[18*(8+1)-1:18*8]));
BIAS #(.value(18'b000001101010011100)) U9  (.q(q[18*(9+1)-1:18*9]));
BIAS #(.value(18'b000000111110000100)) U10 (.q(q[18*(10+1)-1:18*10]));
BIAS #(.value(18'b111111010010010000)) U11 (.q(q[18*(11+1)-1:18*11]));
BIAS #(.value(18'b111110001111010100)) U12 (.q(q[18*(12+1)-1:18*12]));
BIAS #(.value(18'b000011001101100100)) U13 (.q(q[18*(13+1)-1:18*13]));
BIAS #(.value(18'b000000100111001000)) U14 (.q(q[18*(14+1)-1:18*14]));
BIAS #(.value(18'b000001111101011100)) U15 (.q(q[18*(15+1)-1:18*15]));

endmodule