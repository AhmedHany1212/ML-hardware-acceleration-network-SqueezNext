module BIAS_layer1 #(parameter N_adder_tree=64)(q);
output wire [N_adder_tree*18-1:0] q;

BIAS #(.value(18'b111110001101100000)) U0 (.q(q[18*(0+1)-1:18*0])); 
BIAS #(.value(18'b111111010110001100)) U1 (.q(q[18*(1+1)-1:18*1])); 
BIAS #(.value(18'b111111101110111100)) U2 (.q(q[18*(2+1)-1:18*2])); 
BIAS #(.value(18'b000001010011001000)) U3 (.q(q[18*(3+1)-1:18*3])); 
BIAS #(.value(18'b111110001110101100)) U4 (.q(q[18*(4+1)-1:18*4])); 
BIAS #(.value(18'b000000101101001100)) U5 (.q(q[18*(5+1)-1:18*5])); 
BIAS #(.value(18'b000101010110011100)) U6 (.q(q[18*(6+1)-1:18*6])); 
BIAS #(.value(18'b111101111110010000)) U7 (.q(q[18*(7+1)-1:18*7])); 
BIAS #(.value(18'b000001001001010100)) U8 (.q(q[18*(8+1)-1:18*8])); 
BIAS #(.value(18'b111110011010000000)) U9 (.q(q[18*(9+1)-1:18*9])); 
BIAS #(.value(18'b000010001110100100)) U10 (.q(q[18*(10+1)-1:18*10])); 
BIAS #(.value(18'b000000000000010100)) U11 (.q(q[18*(11+1)-1:18*11])); 
BIAS #(.value(18'b111110101000000100)) U12 (.q(q[18*(12+1)-1:18*12])); 
BIAS #(.value(18'b000101101110111000)) U13 (.q(q[18*(13+1)-1:18*13])); 
BIAS #(.value(18'b111111111111010000)) U14 (.q(q[18*(14+1)-1:18*14])); 
BIAS #(.value(18'b111101100101110100)) U15 (.q(q[18*(15+1)-1:18*15])); 
BIAS #(.value(18'b111111000000000000)) U16 (.q(q[18*(16+1)-1:18*16])); 
BIAS #(.value(18'b111111000110101100)) U17 (.q(q[18*(17+1)-1:18*17])); 
BIAS #(.value(18'b000001100100110100)) U18 (.q(q[18*(18+1)-1:18*18])); 
BIAS #(.value(18'b111111010110101100)) U19 (.q(q[18*(19+1)-1:18*19])); 
BIAS #(.value(18'b111100111100101100)) U20 (.q(q[18*(20+1)-1:18*20])); 
BIAS #(.value(18'b000000100110111100)) U21 (.q(q[18*(21+1)-1:18*21])); 
BIAS #(.value(18'b000010011100011000)) U22 (.q(q[18*(22+1)-1:18*22])); 
BIAS #(.value(18'b000000000010101000)) U23 (.q(q[18*(23+1)-1:18*23])); 
BIAS #(.value(18'b000010001010110000)) U24 (.q(q[18*(24+1)-1:18*24])); 
BIAS #(.value(18'b111111110001011000)) U25 (.q(q[18*(25+1)-1:18*25])); 
BIAS #(.value(18'b111111111111011100)) U26 (.q(q[18*(26+1)-1:18*26])); 
BIAS #(.value(18'b000011000001011000)) U27 (.q(q[18*(27+1)-1:18*27])); 
BIAS #(.value(18'b111111000111010100)) U28 (.q(q[18*(28+1)-1:18*28])); 
BIAS #(.value(18'b111111010001110100)) U29 (.q(q[18*(29+1)-1:18*29])); 
BIAS #(.value(18'b000010100001101000)) U30 (.q(q[18*(30+1)-1:18*30])); 
BIAS #(.value(18'b111101110110111100)) U31 (.q(q[18*(31+1)-1:18*31])); 
BIAS #(.value(18'b000010110111000100)) U32 (.q(q[18*(32+1)-1:18*32])); 
BIAS #(.value(18'b000111010010011000)) U33 (.q(q[18*(33+1)-1:18*33])); 
BIAS #(.value(18'b001000010101101100)) U34 (.q(q[18*(34+1)-1:18*34])); 
BIAS #(.value(18'b111111010000010000)) U35 (.q(q[18*(35+1)-1:18*35])); 
BIAS #(.value(18'b111111111111010100)) U36 (.q(q[18*(36+1)-1:18*36])); 
BIAS #(.value(18'b111111010011001000)) U37 (.q(q[18*(37+1)-1:18*37])); 
BIAS #(.value(18'b111110111000010100)) U38 (.q(q[18*(38+1)-1:18*38])); 
BIAS #(.value(18'b111110111010111000)) U39 (.q(q[18*(39+1)-1:18*39])); 
BIAS #(.value(18'b000000000111111100)) U40 (.q(q[18*(40+1)-1:18*40])); 
BIAS #(.value(18'b000001000110011000)) U41 (.q(q[18*(41+1)-1:18*41])); 
BIAS #(.value(18'b111111111100101000)) U42 (.q(q[18*(42+1)-1:18*42])); 
BIAS #(.value(18'b000001101110110000)) U43 (.q(q[18*(43+1)-1:18*43])); 
BIAS #(.value(18'b111111011100101100)) U44 (.q(q[18*(44+1)-1:18*44])); 
BIAS #(.value(18'b000001111000001000)) U45 (.q(q[18*(45+1)-1:18*45])); 
BIAS #(.value(18'b000000001100101000)) U46 (.q(q[18*(46+1)-1:18*46])); 
BIAS #(.value(18'b000111111011000000)) U47 (.q(q[18*(47+1)-1:18*47])); 
BIAS #(.value(18'b111111000011111100)) U48 (.q(q[18*(48+1)-1:18*48])); 
BIAS #(.value(18'b111101110100110000)) U49 (.q(q[18*(49+1)-1:18*49])); 
BIAS #(.value(18'b000010000000011000)) U50 (.q(q[18*(50+1)-1:18*50])); 
BIAS #(.value(18'b111111111111001100)) U51 (.q(q[18*(51+1)-1:18*51])); 
BIAS #(.value(18'b111110000010110000)) U52 (.q(q[18*(52+1)-1:18*52])); 
BIAS #(.value(18'b000000011001010000)) U53 (.q(q[18*(53+1)-1:18*53])); 
BIAS #(.value(18'b000011101010110000)) U54 (.q(q[18*(54+1)-1:18*54])); 
BIAS #(.value(18'b111100110001011000)) U55 (.q(q[18*(55+1)-1:18*55])); 
BIAS #(.value(18'b000001111000101000)) U56 (.q(q[18*(56+1)-1:18*56])); 
BIAS #(.value(18'b111110001100000100)) U57 (.q(q[18*(57+1)-1:18*57])); 
BIAS #(.value(18'b111111101010011000)) U58 (.q(q[18*(58+1)-1:18*58])); 
BIAS #(.value(18'b000010010101111000)) U59 (.q(q[18*(59+1)-1:18*59])); 
BIAS #(.value(18'b000101000110100000)) U60 (.q(q[18*(60+1)-1:18*60])); 
BIAS #(.value(18'b111110100110110100)) U61 (.q(q[18*(61+1)-1:18*61])); 
BIAS #(.value(18'b111111101000010000)) U62 (.q(q[18*(62+1)-1:18*62])); 
BIAS #(.value(18'b000001001100111000)) U63 (.q(q[18*(63+1)-1:18*63])); 

endmodule