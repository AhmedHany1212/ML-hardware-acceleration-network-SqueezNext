

module CONV62 #(parameter N=256,parameter weight_addr_WIDTH=5)(weight_out,weight_addr,clk);
input wire [weight_addr_WIDTH-1:0] weight_addr;
input wire clk;
output wire [N*16-1:0] weight_out ;
W_ROM #(.FILENAME("conv62/CONV62_1.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U0 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv62/CONV62_2.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U1 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv62/CONV62_3.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U2 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv62/CONV62_4.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U3 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv62/CONV62_5.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U4 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv62/CONV62_6.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U5 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv62/CONV62_7.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U6 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv62/CONV62_8.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U7 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv62/CONV62_9.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U8 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv62/CONV62_10.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U9 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv62/CONV62_11.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U10 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv62/CONV62_12.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U11 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv62/CONV62_13.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U12 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv62/CONV62_14.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U13 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv62/CONV62_15.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U14 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv62/CONV62_16.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U15 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv62/CONV62_17.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U16 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv62/CONV62_18.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U17 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv62/CONV62_19.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U18 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv62/CONV62_20.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U19 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv62/CONV62_21.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U20 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv62/CONV62_22.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U21 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv62/CONV62_23.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U22 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv62/CONV62_24.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U23 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv62/CONV62_25.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U24 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv62/CONV62_26.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U25 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv62/CONV62_27.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U26 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv62/CONV62_28.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U27 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv62/CONV62_29.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U28 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv62/CONV62_30.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U29 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv62/CONV62_31.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U30 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv62/CONV62_32.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U31 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv62/CONV62_33.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U32 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv62/CONV62_34.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U33 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv62/CONV62_35.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U34 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv62/CONV62_36.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U35 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv62/CONV62_37.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U36 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv62/CONV62_38.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U37 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv62/CONV62_39.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U38 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv62/CONV62_40.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U39 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv62/CONV62_41.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U40 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv62/CONV62_42.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U41 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv62/CONV62_43.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U42 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv62/CONV62_44.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U43 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv62/CONV62_45.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U44 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv62/CONV62_46.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U45 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv62/CONV62_47.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U46 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv62/CONV62_48.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U47 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv62/CONV62_49.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U48 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv62/CONV62_50.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U49 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv62/CONV62_51.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U50 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv62/CONV62_52.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U51 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv62/CONV62_53.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U52 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv62/CONV62_54.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U53 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv62/CONV62_55.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U54 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv62/CONV62_56.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U55 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv62/CONV62_57.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U56 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv62/CONV62_58.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U57 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv62/CONV62_59.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U58 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv62/CONV62_60.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U59 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv62/CONV62_61.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U60 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv62/CONV62_62.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U61 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv62/CONV62_63.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U62 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv62/CONV62_64.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U63 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(63+1)-1:16*63])); 
W_ROM #(.FILENAME("conv62/CONV62_65.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U64 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(64+1)-1:16*64])); 
W_ROM #(.FILENAME("conv62/CONV62_66.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U65 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(65+1)-1:16*65])); 
W_ROM #(.FILENAME("conv62/CONV62_67.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U66 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(66+1)-1:16*66])); 
W_ROM #(.FILENAME("conv62/CONV62_68.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U67 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(67+1)-1:16*67])); 
W_ROM #(.FILENAME("conv62/CONV62_69.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U68 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(68+1)-1:16*68])); 
W_ROM #(.FILENAME("conv62/CONV62_70.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U69 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(69+1)-1:16*69])); 
W_ROM #(.FILENAME("conv62/CONV62_71.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U70 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(70+1)-1:16*70])); 
W_ROM #(.FILENAME("conv62/CONV62_72.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U71 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(71+1)-1:16*71])); 
W_ROM #(.FILENAME("conv62/CONV62_73.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U72 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(72+1)-1:16*72])); 
W_ROM #(.FILENAME("conv62/CONV62_74.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U73 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(73+1)-1:16*73])); 
W_ROM #(.FILENAME("conv62/CONV62_75.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U74 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(74+1)-1:16*74])); 
W_ROM #(.FILENAME("conv62/CONV62_76.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U75 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(75+1)-1:16*75])); 
W_ROM #(.FILENAME("conv62/CONV62_77.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U76 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(76+1)-1:16*76])); 
W_ROM #(.FILENAME("conv62/CONV62_78.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U77 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(77+1)-1:16*77])); 
W_ROM #(.FILENAME("conv62/CONV62_79.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U78 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(78+1)-1:16*78])); 
W_ROM #(.FILENAME("conv62/CONV62_80.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U79 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(79+1)-1:16*79])); 
W_ROM #(.FILENAME("conv62/CONV62_81.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U80 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(80+1)-1:16*80])); 
W_ROM #(.FILENAME("conv62/CONV62_82.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U81 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(81+1)-1:16*81])); 
W_ROM #(.FILENAME("conv62/CONV62_83.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U82 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(82+1)-1:16*82])); 
W_ROM #(.FILENAME("conv62/CONV62_84.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U83 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(83+1)-1:16*83])); 
W_ROM #(.FILENAME("conv62/CONV62_85.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U84 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(84+1)-1:16*84])); 
W_ROM #(.FILENAME("conv62/CONV62_86.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U85 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(85+1)-1:16*85])); 
W_ROM #(.FILENAME("conv62/CONV62_87.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U86 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(86+1)-1:16*86])); 
W_ROM #(.FILENAME("conv62/CONV62_88.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U87 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(87+1)-1:16*87])); 
W_ROM #(.FILENAME("conv62/CONV62_89.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U88 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(88+1)-1:16*88])); 
W_ROM #(.FILENAME("conv62/CONV62_90.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U89 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(89+1)-1:16*89])); 
W_ROM #(.FILENAME("conv62/CONV62_91.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U90 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(90+1)-1:16*90])); 
W_ROM #(.FILENAME("conv62/CONV62_92.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U91 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(91+1)-1:16*91])); 
W_ROM #(.FILENAME("conv62/CONV62_93.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U92 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(92+1)-1:16*92])); 
W_ROM #(.FILENAME("conv62/CONV62_94.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U93 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(93+1)-1:16*93])); 
W_ROM #(.FILENAME("conv62/CONV62_95.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U94 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(94+1)-1:16*94])); 
W_ROM #(.FILENAME("conv62/CONV62_96.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U95 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(95+1)-1:16*95])); 
W_ROM #(.FILENAME("conv62/CONV62_97.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U96 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(96+1)-1:16*96])); 
W_ROM #(.FILENAME("conv62/CONV62_98.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U97 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(97+1)-1:16*97])); 
W_ROM #(.FILENAME("conv62/CONV62_99.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U98 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(98+1)-1:16*98])); 
W_ROM #(.FILENAME("conv62/CONV62_100.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U99 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(99+1)-1:16*99])); 
W_ROM #(.FILENAME("conv62/CONV62_101.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U100 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(100+1)-1:16*100])); 
W_ROM #(.FILENAME("conv62/CONV62_102.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U101 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(101+1)-1:16*101])); 
W_ROM #(.FILENAME("conv62/CONV62_103.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U102 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(102+1)-1:16*102])); 
W_ROM #(.FILENAME("conv62/CONV62_104.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U103 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(103+1)-1:16*103])); 
W_ROM #(.FILENAME("conv62/CONV62_105.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U104 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(104+1)-1:16*104])); 
W_ROM #(.FILENAME("conv62/CONV62_106.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U105 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(105+1)-1:16*105])); 
W_ROM #(.FILENAME("conv62/CONV62_107.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U106 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(106+1)-1:16*106])); 
W_ROM #(.FILENAME("conv62/CONV62_108.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U107 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(107+1)-1:16*107])); 
W_ROM #(.FILENAME("conv62/CONV62_109.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U108 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(108+1)-1:16*108])); 
W_ROM #(.FILENAME("conv62/CONV62_110.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U109 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(109+1)-1:16*109])); 
W_ROM #(.FILENAME("conv62/CONV62_111.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U110 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(110+1)-1:16*110])); 
W_ROM #(.FILENAME("conv62/CONV62_112.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U111 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(111+1)-1:16*111])); 
W_ROM #(.FILENAME("conv62/CONV62_113.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U112 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(112+1)-1:16*112])); 
W_ROM #(.FILENAME("conv62/CONV62_114.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U113 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(113+1)-1:16*113])); 
W_ROM #(.FILENAME("conv62/CONV62_115.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U114 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(114+1)-1:16*114])); 
W_ROM #(.FILENAME("conv62/CONV62_116.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U115 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(115+1)-1:16*115])); 
W_ROM #(.FILENAME("conv62/CONV62_117.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U116 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(116+1)-1:16*116])); 
W_ROM #(.FILENAME("conv62/CONV62_118.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U117 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(117+1)-1:16*117])); 
W_ROM #(.FILENAME("conv62/CONV62_119.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U118 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(118+1)-1:16*118])); 
W_ROM #(.FILENAME("conv62/CONV62_120.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U119 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(119+1)-1:16*119])); 
W_ROM #(.FILENAME("conv62/CONV62_121.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U120 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(120+1)-1:16*120])); 
W_ROM #(.FILENAME("conv62/CONV62_122.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U121 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(121+1)-1:16*121])); 
W_ROM #(.FILENAME("conv62/CONV62_123.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U122 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(122+1)-1:16*122])); 
W_ROM #(.FILENAME("conv62/CONV62_124.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U123 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(123+1)-1:16*123])); 
W_ROM #(.FILENAME("conv62/CONV62_125.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U124 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(124+1)-1:16*124])); 
W_ROM #(.FILENAME("conv62/CONV62_126.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U125 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(125+1)-1:16*125])); 
W_ROM #(.FILENAME("conv62/CONV62_127.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U126 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(126+1)-1:16*126])); 
W_ROM #(.FILENAME("conv62/CONV62_128.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U127 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(127+1)-1:16*127])); 
W_ROM #(.FILENAME("conv62/CONV62_129.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U128 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(128+1)-1:16*128])); 
W_ROM #(.FILENAME("conv62/CONV62_130.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U129 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(129+1)-1:16*129])); 
W_ROM #(.FILENAME("conv62/CONV62_131.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U130 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(130+1)-1:16*130])); 
W_ROM #(.FILENAME("conv62/CONV62_132.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U131 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(131+1)-1:16*131])); 
W_ROM #(.FILENAME("conv62/CONV62_133.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U132 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(132+1)-1:16*132])); 
W_ROM #(.FILENAME("conv62/CONV62_134.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U133 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(133+1)-1:16*133])); 
W_ROM #(.FILENAME("conv62/CONV62_135.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U134 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(134+1)-1:16*134])); 
W_ROM #(.FILENAME("conv62/CONV62_136.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U135 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(135+1)-1:16*135])); 
W_ROM #(.FILENAME("conv62/CONV62_137.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U136 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(136+1)-1:16*136])); 
W_ROM #(.FILENAME("conv62/CONV62_138.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U137 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(137+1)-1:16*137])); 
W_ROM #(.FILENAME("conv62/CONV62_139.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U138 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(138+1)-1:16*138])); 
W_ROM #(.FILENAME("conv62/CONV62_140.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U139 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(139+1)-1:16*139])); 
W_ROM #(.FILENAME("conv62/CONV62_141.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U140 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(140+1)-1:16*140])); 
W_ROM #(.FILENAME("conv62/CONV62_142.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U141 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(141+1)-1:16*141])); 
W_ROM #(.FILENAME("conv62/CONV62_143.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U142 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(142+1)-1:16*142])); 
W_ROM #(.FILENAME("conv62/CONV62_144.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U143 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(143+1)-1:16*143])); 
W_ROM #(.FILENAME("conv62/CONV62_145.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U144 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(144+1)-1:16*144])); 
W_ROM #(.FILENAME("conv62/CONV62_146.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U145 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(145+1)-1:16*145])); 
W_ROM #(.FILENAME("conv62/CONV62_147.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U146 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(146+1)-1:16*146])); 
W_ROM #(.FILENAME("conv62/CONV62_148.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U147 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(147+1)-1:16*147])); 
W_ROM #(.FILENAME("conv62/CONV62_149.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U148 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(148+1)-1:16*148])); 
W_ROM #(.FILENAME("conv62/CONV62_150.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U149 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(149+1)-1:16*149])); 
W_ROM #(.FILENAME("conv62/CONV62_151.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U150 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(150+1)-1:16*150])); 
W_ROM #(.FILENAME("conv62/CONV62_152.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U151 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(151+1)-1:16*151])); 
W_ROM #(.FILENAME("conv62/CONV62_153.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U152 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(152+1)-1:16*152])); 
W_ROM #(.FILENAME("conv62/CONV62_154.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U153 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(153+1)-1:16*153])); 
W_ROM #(.FILENAME("conv62/CONV62_155.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U154 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(154+1)-1:16*154])); 
W_ROM #(.FILENAME("conv62/CONV62_156.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U155 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(155+1)-1:16*155])); 
W_ROM #(.FILENAME("conv62/CONV62_157.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U156 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(156+1)-1:16*156])); 
W_ROM #(.FILENAME("conv62/CONV62_158.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U157 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(157+1)-1:16*157])); 
W_ROM #(.FILENAME("conv62/CONV62_159.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U158 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(158+1)-1:16*158])); 
W_ROM #(.FILENAME("conv62/CONV62_160.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U159 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(159+1)-1:16*159])); 
W_ROM #(.FILENAME("conv62/CONV62_161.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U160 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(160+1)-1:16*160])); 
W_ROM #(.FILENAME("conv62/CONV62_162.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U161 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(161+1)-1:16*161])); 
W_ROM #(.FILENAME("conv62/CONV62_163.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U162 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(162+1)-1:16*162])); 
W_ROM #(.FILENAME("conv62/CONV62_164.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U163 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(163+1)-1:16*163])); 
W_ROM #(.FILENAME("conv62/CONV62_165.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U164 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(164+1)-1:16*164])); 
W_ROM #(.FILENAME("conv62/CONV62_166.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U165 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(165+1)-1:16*165])); 
W_ROM #(.FILENAME("conv62/CONV62_167.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U166 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(166+1)-1:16*166])); 
W_ROM #(.FILENAME("conv62/CONV62_168.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U167 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(167+1)-1:16*167])); 
W_ROM #(.FILENAME("conv62/CONV62_169.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U168 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(168+1)-1:16*168])); 
W_ROM #(.FILENAME("conv62/CONV62_170.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U169 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(169+1)-1:16*169])); 
W_ROM #(.FILENAME("conv62/CONV62_171.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U170 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(170+1)-1:16*170])); 
W_ROM #(.FILENAME("conv62/CONV62_172.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U171 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(171+1)-1:16*171])); 
W_ROM #(.FILENAME("conv62/CONV62_173.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U172 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(172+1)-1:16*172])); 
W_ROM #(.FILENAME("conv62/CONV62_174.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U173 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(173+1)-1:16*173])); 
W_ROM #(.FILENAME("conv62/CONV62_175.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U174 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(174+1)-1:16*174])); 
W_ROM #(.FILENAME("conv62/CONV62_176.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U175 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(175+1)-1:16*175])); 
W_ROM #(.FILENAME("conv62/CONV62_177.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U176 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(176+1)-1:16*176])); 
W_ROM #(.FILENAME("conv62/CONV62_178.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U177 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(177+1)-1:16*177])); 
W_ROM #(.FILENAME("conv62/CONV62_179.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U178 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(178+1)-1:16*178])); 
W_ROM #(.FILENAME("conv62/CONV62_180.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U179 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(179+1)-1:16*179])); 
W_ROM #(.FILENAME("conv62/CONV62_181.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U180 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(180+1)-1:16*180])); 
W_ROM #(.FILENAME("conv62/CONV62_182.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U181 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(181+1)-1:16*181])); 
W_ROM #(.FILENAME("conv62/CONV62_183.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U182 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(182+1)-1:16*182])); 
W_ROM #(.FILENAME("conv62/CONV62_184.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U183 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(183+1)-1:16*183])); 
W_ROM #(.FILENAME("conv62/CONV62_185.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U184 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(184+1)-1:16*184])); 
W_ROM #(.FILENAME("conv62/CONV62_186.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U185 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(185+1)-1:16*185])); 
W_ROM #(.FILENAME("conv62/CONV62_187.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U186 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(186+1)-1:16*186])); 
W_ROM #(.FILENAME("conv62/CONV62_188.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U187 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(187+1)-1:16*187])); 
W_ROM #(.FILENAME("conv62/CONV62_189.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U188 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(188+1)-1:16*188])); 
W_ROM #(.FILENAME("conv62/CONV62_190.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U189 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(189+1)-1:16*189])); 
W_ROM #(.FILENAME("conv62/CONV62_191.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U190 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(190+1)-1:16*190])); 
W_ROM #(.FILENAME("conv62/CONV62_192.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U191 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(191+1)-1:16*191])); 
W_ROM #(.FILENAME("conv62/CONV62_193.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U192 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(192+1)-1:16*192])); 
W_ROM #(.FILENAME("conv62/CONV62_194.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U193 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(193+1)-1:16*193])); 
W_ROM #(.FILENAME("conv62/CONV62_195.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U194 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(194+1)-1:16*194])); 
W_ROM #(.FILENAME("conv62/CONV62_196.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U195 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(195+1)-1:16*195])); 
W_ROM #(.FILENAME("conv62/CONV62_197.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U196 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(196+1)-1:16*196])); 
W_ROM #(.FILENAME("conv62/CONV62_198.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U197 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(197+1)-1:16*197])); 
W_ROM #(.FILENAME("conv62/CONV62_199.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U198 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(198+1)-1:16*198])); 
W_ROM #(.FILENAME("conv62/CONV62_200.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U199 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(199+1)-1:16*199])); 
W_ROM #(.FILENAME("conv62/CONV62_201.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U200 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(200+1)-1:16*200])); 
W_ROM #(.FILENAME("conv62/CONV62_202.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U201 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(201+1)-1:16*201])); 
W_ROM #(.FILENAME("conv62/CONV62_203.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U202 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(202+1)-1:16*202])); 
W_ROM #(.FILENAME("conv62/CONV62_204.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U203 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(203+1)-1:16*203])); 
W_ROM #(.FILENAME("conv62/CONV62_205.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U204 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(204+1)-1:16*204])); 
W_ROM #(.FILENAME("conv62/CONV62_206.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U205 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(205+1)-1:16*205])); 
W_ROM #(.FILENAME("conv62/CONV62_207.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U206 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(206+1)-1:16*206])); 
W_ROM #(.FILENAME("conv62/CONV62_208.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U207 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(207+1)-1:16*207])); 
W_ROM #(.FILENAME("conv62/CONV62_209.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U208 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(208+1)-1:16*208])); 
W_ROM #(.FILENAME("conv62/CONV62_210.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U209 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(209+1)-1:16*209])); 
W_ROM #(.FILENAME("conv62/CONV62_211.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U210 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(210+1)-1:16*210])); 
W_ROM #(.FILENAME("conv62/CONV62_212.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U211 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(211+1)-1:16*211])); 
W_ROM #(.FILENAME("conv62/CONV62_213.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U212 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(212+1)-1:16*212])); 
W_ROM #(.FILENAME("conv62/CONV62_214.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U213 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(213+1)-1:16*213])); 
W_ROM #(.FILENAME("conv62/CONV62_215.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U214 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(214+1)-1:16*214])); 
W_ROM #(.FILENAME("conv62/CONV62_216.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U215 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(215+1)-1:16*215])); 
W_ROM #(.FILENAME("conv62/CONV62_217.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U216 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(216+1)-1:16*216])); 
W_ROM #(.FILENAME("conv62/CONV62_218.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U217 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(217+1)-1:16*217])); 
W_ROM #(.FILENAME("conv62/CONV62_219.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U218 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(218+1)-1:16*218])); 
W_ROM #(.FILENAME("conv62/CONV62_220.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U219 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(219+1)-1:16*219])); 
W_ROM #(.FILENAME("conv62/CONV62_221.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U220 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(220+1)-1:16*220])); 
W_ROM #(.FILENAME("conv62/CONV62_222.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U221 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(221+1)-1:16*221])); 
W_ROM #(.FILENAME("conv62/CONV62_223.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U222 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(222+1)-1:16*222])); 
W_ROM #(.FILENAME("conv62/CONV62_224.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U223 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(223+1)-1:16*223])); 
W_ROM #(.FILENAME("conv62/CONV62_225.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U224 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(224+1)-1:16*224])); 
W_ROM #(.FILENAME("conv62/CONV62_226.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U225 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(225+1)-1:16*225])); 
W_ROM #(.FILENAME("conv62/CONV62_227.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U226 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(226+1)-1:16*226])); 
W_ROM #(.FILENAME("conv62/CONV62_228.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U227 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(227+1)-1:16*227])); 
W_ROM #(.FILENAME("conv62/CONV62_229.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U228 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(228+1)-1:16*228])); 
W_ROM #(.FILENAME("conv62/CONV62_230.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U229 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(229+1)-1:16*229])); 
W_ROM #(.FILENAME("conv62/CONV62_231.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U230 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(230+1)-1:16*230])); 
W_ROM #(.FILENAME("conv62/CONV62_232.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U231 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(231+1)-1:16*231])); 
W_ROM #(.FILENAME("conv62/CONV62_233.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U232 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(232+1)-1:16*232])); 
W_ROM #(.FILENAME("conv62/CONV62_234.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U233 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(233+1)-1:16*233])); 
W_ROM #(.FILENAME("conv62/CONV62_235.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U234 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(234+1)-1:16*234])); 
W_ROM #(.FILENAME("conv62/CONV62_236.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U235 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(235+1)-1:16*235])); 
W_ROM #(.FILENAME("conv62/CONV62_237.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U236 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(236+1)-1:16*236])); 
W_ROM #(.FILENAME("conv62/CONV62_238.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U237 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(237+1)-1:16*237])); 
W_ROM #(.FILENAME("conv62/CONV62_239.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U238 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(238+1)-1:16*238])); 
W_ROM #(.FILENAME("conv62/CONV62_240.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U239 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(239+1)-1:16*239])); 
W_ROM #(.FILENAME("conv62/CONV62_241.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U240 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(240+1)-1:16*240])); 
W_ROM #(.FILENAME("conv62/CONV62_242.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U241 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(241+1)-1:16*241])); 
W_ROM #(.FILENAME("conv62/CONV62_243.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U242 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(242+1)-1:16*242])); 
W_ROM #(.FILENAME("conv62/CONV62_244.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U243 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(243+1)-1:16*243])); 
W_ROM #(.FILENAME("conv62/CONV62_245.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U244 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(244+1)-1:16*244])); 
W_ROM #(.FILENAME("conv62/CONV62_246.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U245 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(245+1)-1:16*245])); 
W_ROM #(.FILENAME("conv62/CONV62_247.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U246 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(246+1)-1:16*246])); 
W_ROM #(.FILENAME("conv62/CONV62_248.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U247 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(247+1)-1:16*247])); 
W_ROM #(.FILENAME("conv62/CONV62_249.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U248 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(248+1)-1:16*248])); 
W_ROM #(.FILENAME("conv62/CONV62_250.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U249 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(249+1)-1:16*249])); 
W_ROM #(.FILENAME("conv62/CONV62_251.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U250 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(250+1)-1:16*250])); 
W_ROM #(.FILENAME("conv62/CONV62_252.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U251 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(251+1)-1:16*251])); 
W_ROM #(.FILENAME("conv62/CONV62_253.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U252 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(252+1)-1:16*252])); 
W_ROM #(.FILENAME("conv62/CONV62_254.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U253 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(253+1)-1:16*253])); 
W_ROM #(.FILENAME("conv62/CONV62_255.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U254 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(254+1)-1:16*254])); 
W_ROM #(.FILENAME("conv62/CONV62_256.txt"),.weight_addr_WIDTH(5),.NO_ROWS(32)) U255 (.clk(clk),.weight_addr(weight_addr),.weight_out(weight_out[16*(255+1)-1:16*255])); 


endmodule
