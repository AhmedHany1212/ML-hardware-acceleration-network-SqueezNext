module CONV17 #(parameter N=256,parameter ADDR_WIDTH=4)(addr,clk,q);
input wire [ADDR_WIDTH-1:0] addr;
output wire [N*16-1:0] q ;
input clk;
W_ROM#(.FILENAME("conv17/CONV17_1.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U0 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(0+1)-1:16*0])); 
W_ROM#(.FILENAME("conv17/CONV17_2.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U1 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(1+1)-1:16*1])); 
W_ROM#(.FILENAME("conv17/CONV17_3.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U2 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(2+1)-1:16*2])); 
W_ROM#(.FILENAME("conv17/CONV17_4.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U3 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(3+1)-1:16*3])); 
W_ROM#(.FILENAME("conv17/CONV17_5.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U4 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(4+1)-1:16*4])); 
W_ROM#(.FILENAME("conv17/CONV17_6.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U5 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(5+1)-1:16*5])); 
W_ROM#(.FILENAME("conv17/CONV17_7.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U6 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(6+1)-1:16*6])); 
W_ROM#(.FILENAME("conv17/CONV17_8.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U7 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(7+1)-1:16*7])); 
W_ROM#(.FILENAME("conv17/CONV17_9.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U8 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(8+1)-1:16*8])); 
W_ROM#(.FILENAME("conv17/CONV17_10.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U9 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(9+1)-1:16*9])); 
W_ROM#(.FILENAME("conv17/CONV17_11.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U10 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(10+1)-1:16*10])); 
W_ROM#(.FILENAME("conv17/CONV17_12.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U11 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(11+1)-1:16*11])); 
W_ROM#(.FILENAME("conv17/CONV17_13.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U12 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(12+1)-1:16*12])); 
W_ROM#(.FILENAME("conv17/CONV17_14.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U13 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(13+1)-1:16*13])); 
W_ROM#(.FILENAME("conv17/CONV17_15.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U14 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(14+1)-1:16*14])); 
W_ROM#(.FILENAME("conv17/CONV17_16.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U15 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(15+1)-1:16*15])); 
W_ROM#(.FILENAME("conv17/CONV17_17.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U16 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(16+1)-1:16*16])); 
W_ROM#(.FILENAME("conv17/CONV17_18.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U17 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(17+1)-1:16*17])); 
W_ROM#(.FILENAME("conv17/CONV17_19.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U18 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(18+1)-1:16*18])); 
W_ROM#(.FILENAME("conv17/CONV17_20.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U19 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(19+1)-1:16*19])); 
W_ROM#(.FILENAME("conv17/CONV17_21.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U20 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(20+1)-1:16*20])); 
W_ROM#(.FILENAME("conv17/CONV17_22.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U21 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(21+1)-1:16*21])); 
W_ROM#(.FILENAME("conv17/CONV17_23.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U22 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(22+1)-1:16*22])); 
W_ROM#(.FILENAME("conv17/CONV17_24.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U23 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(23+1)-1:16*23])); 
W_ROM#(.FILENAME("conv17/CONV17_25.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U24 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(24+1)-1:16*24])); 
W_ROM#(.FILENAME("conv17/CONV17_26.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U25 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(25+1)-1:16*25])); 
W_ROM#(.FILENAME("conv17/CONV17_27.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U26 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(26+1)-1:16*26])); 
W_ROM#(.FILENAME("conv17/CONV17_28.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U27 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(27+1)-1:16*27])); 
W_ROM#(.FILENAME("conv17/CONV17_29.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U28 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(28+1)-1:16*28])); 
W_ROM#(.FILENAME("conv17/CONV17_30.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U29 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(29+1)-1:16*29])); 
W_ROM#(.FILENAME("conv17/CONV17_31.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U30 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(30+1)-1:16*30])); 
W_ROM#(.FILENAME("conv17/CONV17_32.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U31 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(31+1)-1:16*31])); 
W_ROM#(.FILENAME("conv17/CONV17_33.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U32 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(32+1)-1:16*32])); 
W_ROM#(.FILENAME("conv17/CONV17_34.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U33 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(33+1)-1:16*33])); 
W_ROM#(.FILENAME("conv17/CONV17_35.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U34 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(34+1)-1:16*34])); 
W_ROM#(.FILENAME("conv17/CONV17_36.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U35 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(35+1)-1:16*35])); 
W_ROM#(.FILENAME("conv17/CONV17_37.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U36 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(36+1)-1:16*36])); 
W_ROM#(.FILENAME("conv17/CONV17_38.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U37 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(37+1)-1:16*37])); 
W_ROM#(.FILENAME("conv17/CONV17_39.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U38 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(38+1)-1:16*38])); 
W_ROM#(.FILENAME("conv17/CONV17_40.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U39 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(39+1)-1:16*39])); 
W_ROM#(.FILENAME("conv17/CONV17_41.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U40 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(40+1)-1:16*40])); 
W_ROM#(.FILENAME("conv17/CONV17_42.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U41 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(41+1)-1:16*41])); 
W_ROM#(.FILENAME("conv17/CONV17_43.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U42 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(42+1)-1:16*42])); 
W_ROM#(.FILENAME("conv17/CONV17_44.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U43 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(43+1)-1:16*43])); 
W_ROM#(.FILENAME("conv17/CONV17_45.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U44 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(44+1)-1:16*44])); 
W_ROM#(.FILENAME("conv17/CONV17_46.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U45 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(45+1)-1:16*45])); 
W_ROM#(.FILENAME("conv17/CONV17_47.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U46 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(46+1)-1:16*46])); 
W_ROM#(.FILENAME("conv17/CONV17_48.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U47 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(47+1)-1:16*47])); 
W_ROM#(.FILENAME("conv17/CONV17_49.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U48 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(48+1)-1:16*48])); 
W_ROM#(.FILENAME("conv17/CONV17_50.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U49 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(49+1)-1:16*49])); 
W_ROM#(.FILENAME("conv17/CONV17_51.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U50 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(50+1)-1:16*50])); 
W_ROM#(.FILENAME("conv17/CONV17_52.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U51 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(51+1)-1:16*51])); 
W_ROM#(.FILENAME("conv17/CONV17_53.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U52 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(52+1)-1:16*52])); 
W_ROM#(.FILENAME("conv17/CONV17_54.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U53 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(53+1)-1:16*53])); 
W_ROM#(.FILENAME("conv17/CONV17_55.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U54 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(54+1)-1:16*54])); 
W_ROM#(.FILENAME("conv17/CONV17_56.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U55 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(55+1)-1:16*55])); 
W_ROM#(.FILENAME("conv17/CONV17_57.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U56 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(56+1)-1:16*56])); 
W_ROM#(.FILENAME("conv17/CONV17_58.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U57 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(57+1)-1:16*57])); 
W_ROM#(.FILENAME("conv17/CONV17_59.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U58 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(58+1)-1:16*58])); 
W_ROM#(.FILENAME("conv17/CONV17_60.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U59 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(59+1)-1:16*59])); 
W_ROM#(.FILENAME("conv17/CONV17_61.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U60 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(60+1)-1:16*60])); 
W_ROM#(.FILENAME("conv17/CONV17_62.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U61 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(61+1)-1:16*61])); 
W_ROM#(.FILENAME("conv17/CONV17_63.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U62 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(62+1)-1:16*62])); 
W_ROM#(.FILENAME("conv17/CONV17_64.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U63 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(63+1)-1:16*63])); 
W_ROM#(.FILENAME("conv17/CONV17_65.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U64 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(64+1)-1:16*64])); 
W_ROM#(.FILENAME("conv17/CONV17_66.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U65 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(65+1)-1:16*65])); 
W_ROM#(.FILENAME("conv17/CONV17_67.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U66 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(66+1)-1:16*66])); 
W_ROM#(.FILENAME("conv17/CONV17_68.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U67 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(67+1)-1:16*67])); 
W_ROM#(.FILENAME("conv17/CONV17_69.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U68 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(68+1)-1:16*68])); 
W_ROM#(.FILENAME("conv17/CONV17_70.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U69 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(69+1)-1:16*69])); 
W_ROM#(.FILENAME("conv17/CONV17_71.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U70 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(70+1)-1:16*70])); 
W_ROM#(.FILENAME("conv17/CONV17_72.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U71 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(71+1)-1:16*71])); 
W_ROM#(.FILENAME("conv17/CONV17_73.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U72 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(72+1)-1:16*72])); 
W_ROM#(.FILENAME("conv17/CONV17_74.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U73 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(73+1)-1:16*73])); 
W_ROM#(.FILENAME("conv17/CONV17_75.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U74 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(74+1)-1:16*74])); 
W_ROM#(.FILENAME("conv17/CONV17_76.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U75 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(75+1)-1:16*75])); 
W_ROM#(.FILENAME("conv17/CONV17_77.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U76 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(76+1)-1:16*76])); 
W_ROM#(.FILENAME("conv17/CONV17_78.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U77 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(77+1)-1:16*77])); 
W_ROM#(.FILENAME("conv17/CONV17_79.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U78 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(78+1)-1:16*78])); 
W_ROM#(.FILENAME("conv17/CONV17_80.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U79 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(79+1)-1:16*79])); 
W_ROM#(.FILENAME("conv17/CONV17_81.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U80 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(80+1)-1:16*80])); 
W_ROM#(.FILENAME("conv17/CONV17_82.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U81 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(81+1)-1:16*81])); 
W_ROM#(.FILENAME("conv17/CONV17_83.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U82 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(82+1)-1:16*82])); 
W_ROM#(.FILENAME("conv17/CONV17_84.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U83 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(83+1)-1:16*83])); 
W_ROM#(.FILENAME("conv17/CONV17_85.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U84 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(84+1)-1:16*84])); 
W_ROM#(.FILENAME("conv17/CONV17_86.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U85 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(85+1)-1:16*85])); 
W_ROM#(.FILENAME("conv17/CONV17_87.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U86 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(86+1)-1:16*86])); 
W_ROM#(.FILENAME("conv17/CONV17_88.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U87 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(87+1)-1:16*87])); 
W_ROM#(.FILENAME("conv17/CONV17_89.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U88 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(88+1)-1:16*88])); 
W_ROM#(.FILENAME("conv17/CONV17_90.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U89 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(89+1)-1:16*89])); 
W_ROM#(.FILENAME("conv17/CONV17_91.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U90 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(90+1)-1:16*90])); 
W_ROM#(.FILENAME("conv17/CONV17_92.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U91 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(91+1)-1:16*91])); 
W_ROM#(.FILENAME("conv17/CONV17_93.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U92 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(92+1)-1:16*92])); 
W_ROM#(.FILENAME("conv17/CONV17_94.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U93 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(93+1)-1:16*93])); 
W_ROM#(.FILENAME("conv17/CONV17_95.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U94 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(94+1)-1:16*94])); 
W_ROM#(.FILENAME("conv17/CONV17_96.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U95 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(95+1)-1:16*95])); 
W_ROM#(.FILENAME("conv17/CONV17_97.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U96 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(96+1)-1:16*96])); 
W_ROM#(.FILENAME("conv17/CONV17_98.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U97 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(97+1)-1:16*97])); 
W_ROM#(.FILENAME("conv17/CONV17_99.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U98 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(98+1)-1:16*98])); 
W_ROM#(.FILENAME("conv17/CONV17_100.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U99 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(99+1)-1:16*99])); 
W_ROM#(.FILENAME("conv17/CONV17_101.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U100 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(100+1)-1:16*100])); 
W_ROM#(.FILENAME("conv17/CONV17_102.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U101 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(101+1)-1:16*101])); 
W_ROM#(.FILENAME("conv17/CONV17_103.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U102 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(102+1)-1:16*102])); 
W_ROM#(.FILENAME("conv17/CONV17_104.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U103 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(103+1)-1:16*103])); 
W_ROM#(.FILENAME("conv17/CONV17_105.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U104 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(104+1)-1:16*104])); 
W_ROM#(.FILENAME("conv17/CONV17_106.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U105 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(105+1)-1:16*105])); 
W_ROM#(.FILENAME("conv17/CONV17_107.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U106 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(106+1)-1:16*106])); 
W_ROM#(.FILENAME("conv17/CONV17_108.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U107 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(107+1)-1:16*107])); 
W_ROM#(.FILENAME("conv17/CONV17_109.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U108 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(108+1)-1:16*108])); 
W_ROM#(.FILENAME("conv17/CONV17_110.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U109 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(109+1)-1:16*109])); 
W_ROM#(.FILENAME("conv17/CONV17_111.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U110 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(110+1)-1:16*110])); 
W_ROM#(.FILENAME("conv17/CONV17_112.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U111 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(111+1)-1:16*111])); 
W_ROM#(.FILENAME("conv17/CONV17_113.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U112 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(112+1)-1:16*112])); 
W_ROM#(.FILENAME("conv17/CONV17_114.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U113 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(113+1)-1:16*113])); 
W_ROM#(.FILENAME("conv17/CONV17_115.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U114 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(114+1)-1:16*114])); 
W_ROM#(.FILENAME("conv17/CONV17_116.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U115 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(115+1)-1:16*115])); 
W_ROM#(.FILENAME("conv17/CONV17_117.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U116 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(116+1)-1:16*116])); 
W_ROM#(.FILENAME("conv17/CONV17_118.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U117 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(117+1)-1:16*117])); 
W_ROM#(.FILENAME("conv17/CONV17_119.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U118 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(118+1)-1:16*118])); 
W_ROM#(.FILENAME("conv17/CONV17_120.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U119 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(119+1)-1:16*119])); 
W_ROM#(.FILENAME("conv17/CONV17_121.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U120 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(120+1)-1:16*120])); 
W_ROM#(.FILENAME("conv17/CONV17_122.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U121 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(121+1)-1:16*121])); 
W_ROM#(.FILENAME("conv17/CONV17_123.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U122 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(122+1)-1:16*122])); 
W_ROM#(.FILENAME("conv17/CONV17_124.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U123 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(123+1)-1:16*123])); 
W_ROM#(.FILENAME("conv17/CONV17_125.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U124 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(124+1)-1:16*124])); 
W_ROM#(.FILENAME("conv17/CONV17_126.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U125 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(125+1)-1:16*125])); 
W_ROM#(.FILENAME("conv17/CONV17_127.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U126 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(126+1)-1:16*126])); 
W_ROM#(.FILENAME("conv17/CONV17_128.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U127 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(127+1)-1:16*127])); 
W_ROM#(.FILENAME("conv17/CONV17_129.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U128 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(128+1)-1:16*128])); 
W_ROM#(.FILENAME("conv17/CONV17_130.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U129 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(129+1)-1:16*129])); 
W_ROM#(.FILENAME("conv17/CONV17_131.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U130 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(130+1)-1:16*130])); 
W_ROM#(.FILENAME("conv17/CONV17_132.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U131 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(131+1)-1:16*131])); 
W_ROM#(.FILENAME("conv17/CONV17_133.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U132 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(132+1)-1:16*132])); 
W_ROM#(.FILENAME("conv17/CONV17_134.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U133 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(133+1)-1:16*133])); 
W_ROM#(.FILENAME("conv17/CONV17_135.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U134 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(134+1)-1:16*134])); 
W_ROM#(.FILENAME("conv17/CONV17_136.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U135 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(135+1)-1:16*135])); 
W_ROM#(.FILENAME("conv17/CONV17_137.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U136 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(136+1)-1:16*136])); 
W_ROM#(.FILENAME("conv17/CONV17_138.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U137 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(137+1)-1:16*137])); 
W_ROM#(.FILENAME("conv17/CONV17_139.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U138 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(138+1)-1:16*138])); 
W_ROM#(.FILENAME("conv17/CONV17_140.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U139 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(139+1)-1:16*139])); 
W_ROM#(.FILENAME("conv17/CONV17_141.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U140 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(140+1)-1:16*140])); 
W_ROM#(.FILENAME("conv17/CONV17_142.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U141 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(141+1)-1:16*141])); 
W_ROM#(.FILENAME("conv17/CONV17_143.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U142 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(142+1)-1:16*142])); 
W_ROM#(.FILENAME("conv17/CONV17_144.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U143 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(143+1)-1:16*143])); 
W_ROM#(.FILENAME("conv17/CONV17_145.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U144 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(144+1)-1:16*144])); 
W_ROM#(.FILENAME("conv17/CONV17_146.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U145 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(145+1)-1:16*145])); 
W_ROM#(.FILENAME("conv17/CONV17_147.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U146 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(146+1)-1:16*146])); 
W_ROM#(.FILENAME("conv17/CONV17_148.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U147 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(147+1)-1:16*147])); 
W_ROM#(.FILENAME("conv17/CONV17_149.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U148 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(148+1)-1:16*148])); 
W_ROM#(.FILENAME("conv17/CONV17_150.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U149 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(149+1)-1:16*149])); 
W_ROM#(.FILENAME("conv17/CONV17_151.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U150 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(150+1)-1:16*150])); 
W_ROM#(.FILENAME("conv17/CONV17_152.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U151 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(151+1)-1:16*151])); 
W_ROM#(.FILENAME("conv17/CONV17_153.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U152 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(152+1)-1:16*152])); 
W_ROM#(.FILENAME("conv17/CONV17_154.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U153 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(153+1)-1:16*153])); 
W_ROM#(.FILENAME("conv17/CONV17_155.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U154 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(154+1)-1:16*154])); 
W_ROM#(.FILENAME("conv17/CONV17_156.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U155 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(155+1)-1:16*155])); 
W_ROM#(.FILENAME("conv17/CONV17_157.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U156 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(156+1)-1:16*156])); 
W_ROM#(.FILENAME("conv17/CONV17_158.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U157 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(157+1)-1:16*157])); 
W_ROM#(.FILENAME("conv17/CONV17_159.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U158 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(158+1)-1:16*158])); 
W_ROM#(.FILENAME("conv17/CONV17_160.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U159 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(159+1)-1:16*159])); 
W_ROM#(.FILENAME("conv17/CONV17_161.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U160 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(160+1)-1:16*160])); 
W_ROM#(.FILENAME("conv17/CONV17_162.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U161 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(161+1)-1:16*161])); 
W_ROM#(.FILENAME("conv17/CONV17_163.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U162 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(162+1)-1:16*162])); 
W_ROM#(.FILENAME("conv17/CONV17_164.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U163 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(163+1)-1:16*163])); 
W_ROM#(.FILENAME("conv17/CONV17_165.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U164 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(164+1)-1:16*164])); 
W_ROM#(.FILENAME("conv17/CONV17_166.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U165 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(165+1)-1:16*165])); 
W_ROM#(.FILENAME("conv17/CONV17_167.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U166 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(166+1)-1:16*166])); 
W_ROM#(.FILENAME("conv17/CONV17_168.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U167 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(167+1)-1:16*167])); 
W_ROM#(.FILENAME("conv17/CONV17_169.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U168 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(168+1)-1:16*168])); 
W_ROM#(.FILENAME("conv17/CONV17_170.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U169 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(169+1)-1:16*169])); 
W_ROM#(.FILENAME("conv17/CONV17_171.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U170 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(170+1)-1:16*170])); 
W_ROM#(.FILENAME("conv17/CONV17_172.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U171 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(171+1)-1:16*171])); 
W_ROM#(.FILENAME("conv17/CONV17_173.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U172 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(172+1)-1:16*172])); 
W_ROM#(.FILENAME("conv17/CONV17_174.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U173 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(173+1)-1:16*173])); 
W_ROM#(.FILENAME("conv17/CONV17_175.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U174 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(174+1)-1:16*174])); 
W_ROM#(.FILENAME("conv17/CONV17_176.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U175 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(175+1)-1:16*175])); 
W_ROM#(.FILENAME("conv17/CONV17_177.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U176 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(176+1)-1:16*176])); 
W_ROM#(.FILENAME("conv17/CONV17_178.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U177 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(177+1)-1:16*177])); 
W_ROM#(.FILENAME("conv17/CONV17_179.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U178 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(178+1)-1:16*178])); 
W_ROM#(.FILENAME("conv17/CONV17_180.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U179 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(179+1)-1:16*179])); 
W_ROM#(.FILENAME("conv17/CONV17_181.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U180 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(180+1)-1:16*180])); 
W_ROM#(.FILENAME("conv17/CONV17_182.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U181 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(181+1)-1:16*181])); 
W_ROM#(.FILENAME("conv17/CONV17_183.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U182 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(182+1)-1:16*182])); 
W_ROM#(.FILENAME("conv17/CONV17_184.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U183 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(183+1)-1:16*183])); 
W_ROM#(.FILENAME("conv17/CONV17_185.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U184 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(184+1)-1:16*184])); 
W_ROM#(.FILENAME("conv17/CONV17_186.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U185 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(185+1)-1:16*185])); 
W_ROM#(.FILENAME("conv17/CONV17_187.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U186 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(186+1)-1:16*186])); 
W_ROM#(.FILENAME("conv17/CONV17_188.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U187 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(187+1)-1:16*187])); 
W_ROM#(.FILENAME("conv17/CONV17_189.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U188 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(188+1)-1:16*188])); 
W_ROM#(.FILENAME("conv17/CONV17_190.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U189 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(189+1)-1:16*189])); 
W_ROM#(.FILENAME("conv17/CONV17_191.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U190 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(190+1)-1:16*190])); 
W_ROM#(.FILENAME("conv17/CONV17_192.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U191 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(191+1)-1:16*191])); 
W_ROM#(.FILENAME("conv17/CONV17_193.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U192 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(192+1)-1:16*192])); 
W_ROM#(.FILENAME("conv17/CONV17_194.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U193 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(193+1)-1:16*193])); 
W_ROM#(.FILENAME("conv17/CONV17_195.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U194 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(194+1)-1:16*194])); 
W_ROM#(.FILENAME("conv17/CONV17_196.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U195 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(195+1)-1:16*195])); 
W_ROM#(.FILENAME("conv17/CONV17_197.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U196 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(196+1)-1:16*196])); 
W_ROM#(.FILENAME("conv17/CONV17_198.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U197 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(197+1)-1:16*197])); 
W_ROM#(.FILENAME("conv17/CONV17_199.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U198 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(198+1)-1:16*198])); 
W_ROM#(.FILENAME("conv17/CONV17_200.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U199 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(199+1)-1:16*199])); 
W_ROM#(.FILENAME("conv17/CONV17_201.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U200 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(200+1)-1:16*200])); 
W_ROM#(.FILENAME("conv17/CONV17_202.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U201 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(201+1)-1:16*201])); 
W_ROM#(.FILENAME("conv17/CONV17_203.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U202 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(202+1)-1:16*202])); 
W_ROM#(.FILENAME("conv17/CONV17_204.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U203 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(203+1)-1:16*203])); 
W_ROM#(.FILENAME("conv17/CONV17_205.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U204 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(204+1)-1:16*204])); 
W_ROM#(.FILENAME("conv17/CONV17_206.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U205 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(205+1)-1:16*205])); 
W_ROM#(.FILENAME("conv17/CONV17_207.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U206 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(206+1)-1:16*206])); 
W_ROM#(.FILENAME("conv17/CONV17_208.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U207 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(207+1)-1:16*207])); 
W_ROM#(.FILENAME("conv17/CONV17_209.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U208 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(208+1)-1:16*208])); 
W_ROM#(.FILENAME("conv17/CONV17_210.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U209 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(209+1)-1:16*209])); 
W_ROM#(.FILENAME("conv17/CONV17_211.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U210 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(210+1)-1:16*210])); 
W_ROM#(.FILENAME("conv17/CONV17_212.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U211 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(211+1)-1:16*211])); 
W_ROM#(.FILENAME("conv17/CONV17_213.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U212 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(212+1)-1:16*212])); 
W_ROM#(.FILENAME("conv17/CONV17_214.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U213 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(213+1)-1:16*213])); 
W_ROM#(.FILENAME("conv17/CONV17_215.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U214 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(214+1)-1:16*214])); 
W_ROM#(.FILENAME("conv17/CONV17_216.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U215 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(215+1)-1:16*215])); 
W_ROM#(.FILENAME("conv17/CONV17_217.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U216 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(216+1)-1:16*216])); 
W_ROM#(.FILENAME("conv17/CONV17_218.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U217 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(217+1)-1:16*217])); 
W_ROM#(.FILENAME("conv17/CONV17_219.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U218 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(218+1)-1:16*218])); 
W_ROM#(.FILENAME("conv17/CONV17_220.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U219 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(219+1)-1:16*219])); 
W_ROM#(.FILENAME("conv17/CONV17_221.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U220 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(220+1)-1:16*220])); 
W_ROM#(.FILENAME("conv17/CONV17_222.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U221 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(221+1)-1:16*221])); 
W_ROM#(.FILENAME("conv17/CONV17_223.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U222 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(222+1)-1:16*222])); 
W_ROM#(.FILENAME("conv17/CONV17_224.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U223 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(223+1)-1:16*223])); 
W_ROM#(.FILENAME("conv17/CONV17_225.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U224 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(224+1)-1:16*224])); 
W_ROM#(.FILENAME("conv17/CONV17_226.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U225 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(225+1)-1:16*225])); 
W_ROM#(.FILENAME("conv17/CONV17_227.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U226 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(226+1)-1:16*226])); 
W_ROM#(.FILENAME("conv17/CONV17_228.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U227 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(227+1)-1:16*227])); 
W_ROM#(.FILENAME("conv17/CONV17_229.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U228 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(228+1)-1:16*228])); 
W_ROM#(.FILENAME("conv17/CONV17_230.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U229 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(229+1)-1:16*229])); 
W_ROM#(.FILENAME("conv17/CONV17_231.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U230 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(230+1)-1:16*230])); 
W_ROM#(.FILENAME("conv17/CONV17_232.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U231 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(231+1)-1:16*231])); 
W_ROM#(.FILENAME("conv17/CONV17_233.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U232 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(232+1)-1:16*232])); 
W_ROM#(.FILENAME("conv17/CONV17_234.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U233 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(233+1)-1:16*233])); 
W_ROM#(.FILENAME("conv17/CONV17_235.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U234 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(234+1)-1:16*234])); 
W_ROM#(.FILENAME("conv17/CONV17_236.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U235 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(235+1)-1:16*235])); 
W_ROM#(.FILENAME("conv17/CONV17_237.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U236 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(236+1)-1:16*236])); 
W_ROM#(.FILENAME("conv17/CONV17_238.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U237 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(237+1)-1:16*237])); 
W_ROM#(.FILENAME("conv17/CONV17_239.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U238 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(238+1)-1:16*238])); 
W_ROM#(.FILENAME("conv17/CONV17_240.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U239 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(239+1)-1:16*239])); 
W_ROM#(.FILENAME("conv17/CONV17_241.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U240 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(240+1)-1:16*240])); 
W_ROM#(.FILENAME("conv17/CONV17_242.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U241 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(241+1)-1:16*241])); 
W_ROM#(.FILENAME("conv17/CONV17_243.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U242 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(242+1)-1:16*242])); 
W_ROM#(.FILENAME("conv17/CONV17_244.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U243 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(243+1)-1:16*243])); 
W_ROM#(.FILENAME("conv17/CONV17_245.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U244 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(244+1)-1:16*244])); 
W_ROM#(.FILENAME("conv17/CONV17_246.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U245 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(245+1)-1:16*245])); 
W_ROM#(.FILENAME("conv17/CONV17_247.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U246 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(246+1)-1:16*246])); 
W_ROM#(.FILENAME("conv17/CONV17_248.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U247 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(247+1)-1:16*247])); 
W_ROM#(.FILENAME("conv17/CONV17_249.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U248 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(248+1)-1:16*248])); 
W_ROM#(.FILENAME("conv17/CONV17_250.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U249 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(249+1)-1:16*249])); 
W_ROM#(.FILENAME("conv17/CONV17_251.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U250 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(250+1)-1:16*250])); 
W_ROM#(.FILENAME("conv17/CONV17_252.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U251 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(251+1)-1:16*251])); 
W_ROM#(.FILENAME("conv17/CONV17_253.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U252 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(252+1)-1:16*252])); 
W_ROM#(.FILENAME("conv17/CONV17_254.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U253 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(253+1)-1:16*253])); 
W_ROM#(.FILENAME("conv17/CONV17_255.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U254 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(254+1)-1:16*254])); 
W_ROM#(.FILENAME("conv17/CONV17_256.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U255 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(255+1)-1:16*255])); 


endmodule
