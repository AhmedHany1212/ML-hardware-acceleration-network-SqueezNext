module CONV5 #(parameter N=32,parameter weight_addr_WIDTH=4)(addr,clk,q);
input wire [weight_addr_WIDTH-1:0] addr;
input wire clk;
output wire [N*16-1:0] q ;
W_ROM #(.FILENAME("CONV5/CONV5_1.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U0 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("CONV5/CONV5_2.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U1 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("CONV5/CONV5_3.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U2 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("CONV5/CONV5_4.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U3 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("CONV5/CONV5_5.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U4 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("CONV5/CONV5_6.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U5 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("CONV5/CONV5_7.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U6 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("CONV5/CONV5_8.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U7 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("CONV5/CONV5_9.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U8 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("CONV5/CONV5_10.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U9 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("CONV5/CONV5_11.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U10 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("CONV5/CONV5_12.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U11 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("CONV5/CONV5_13.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U12 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("CONV5/CONV5_14.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U13 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("CONV5/CONV5_15.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U14 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("CONV5/CONV5_16.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U15 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("CONV5/CONV5_17.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U16 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("CONV5/CONV5_18.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U17 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("CONV5/CONV5_19.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U18 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("CONV5/CONV5_20.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U19 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("CONV5/CONV5_21.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U20 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("CONV5/CONV5_22.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U21 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("CONV5/CONV5_23.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U22 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("CONV5/CONV5_24.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U23 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("CONV5/CONV5_25.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U24 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("CONV5/CONV5_26.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U25 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("CONV5/CONV5_27.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U26 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("CONV5/CONV5_28.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U27 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("CONV5/CONV5_29.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U28 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("CONV5/CONV5_30.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U29 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("CONV5/CONV5_31.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U30 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("CONV5/CONV5_32.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U31 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(31+1)-1:16*31])); 


endmodule