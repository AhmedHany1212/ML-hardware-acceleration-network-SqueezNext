module CONV3 #(parameter N=128,parameter weight_addr_WIDTH=3)(weight_addr,clk,weight_out);
input wire [weight_addr_WIDTH-1:0] weight_addr;
output wire [N*16-1:0] weight_out ;
input clk;
W_ROM #(.FILENAME("conv3/CONV3_1.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U0 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv3/CONV3_2.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U1 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(1+1)-1:16*1])); 
W_ROM#(.FILENAME("conv3/CONV3_3.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U2 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(2+1)-1:16*2])); 
W_ROM#(.FILENAME("conv3/CONV3_4.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U3 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(3+1)-1:16*3])); 
W_ROM#(.FILENAME("conv3/CONV3_5.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U4 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(4+1)-1:16*4])); 
W_ROM#(.FILENAME("conv3/CONV3_6.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U5 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(5+1)-1:16*5])); 
W_ROM#(.FILENAME("conv3/CONV3_7.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U6 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(6+1)-1:16*6])); 
W_ROM#(.FILENAME("conv3/CONV3_8.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U7 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(7+1)-1:16*7])); 
W_ROM#(.FILENAME("conv3/CONV3_9.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U8 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(8+1)-1:16*8])); 
W_ROM#(.FILENAME("conv3/CONV3_10.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U9 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(9+1)-1:16*9])); 
W_ROM#(.FILENAME("conv3/CONV3_11.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U10 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(10+1)-1:16*10])); 
W_ROM#(.FILENAME("conv3/CONV3_12.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U11 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(11+1)-1:16*11])); 
W_ROM#(.FILENAME("conv3/CONV3_13.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U12 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(12+1)-1:16*12])); 
W_ROM#(.FILENAME("conv3/CONV3_14.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U13 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(13+1)-1:16*13])); 
W_ROM#(.FILENAME("conv3/CONV3_15.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U14 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(14+1)-1:16*14])); 
W_ROM#(.FILENAME("conv3/CONV3_16.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U15 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(15+1)-1:16*15])); 
W_ROM#(.FILENAME("conv3/CONV3_17.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U16 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(16+1)-1:16*16])); 
W_ROM#(.FILENAME("conv3/CONV3_18.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U17 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(17+1)-1:16*17])); 
W_ROM#(.FILENAME("conv3/CONV3_19.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U18 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(18+1)-1:16*18])); 
W_ROM#(.FILENAME("conv3/CONV3_20.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U19 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(19+1)-1:16*19])); 
W_ROM#(.FILENAME("conv3/CONV3_21.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U20 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(20+1)-1:16*20])); 
W_ROM#(.FILENAME("conv3/CONV3_22.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U21 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(21+1)-1:16*21])); 
W_ROM#(.FILENAME("conv3/CONV3_23.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U22 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(22+1)-1:16*22])); 
W_ROM#(.FILENAME("conv3/CONV3_24.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U23 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(23+1)-1:16*23])); 
W_ROM#(.FILENAME("conv3/CONV3_25.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U24 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(24+1)-1:16*24])); 
W_ROM#(.FILENAME("conv3/CONV3_26.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U25 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(25+1)-1:16*25])); 
W_ROM#(.FILENAME("conv3/CONV3_27.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U26 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(26+1)-1:16*26])); 
W_ROM#(.FILENAME("conv3/CONV3_28.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U27 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(27+1)-1:16*27])); 
W_ROM#(.FILENAME("conv3/CONV3_29.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U28 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(28+1)-1:16*28])); 
W_ROM#(.FILENAME("conv3/CONV3_30.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U29 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(29+1)-1:16*29])); 
W_ROM#(.FILENAME("conv3/CONV3_31.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U30 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(30+1)-1:16*30])); 
W_ROM#(.FILENAME("conv3/CONV3_32.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U31 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(31+1)-1:16*31])); 
W_ROM#(.FILENAME("conv3/CONV3_33.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U32 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(32+1)-1:16*32])); 
W_ROM#(.FILENAME("conv3/CONV3_34.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U33 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(33+1)-1:16*33])); 
W_ROM#(.FILENAME("conv3/CONV3_35.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U34 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(34+1)-1:16*34])); 
W_ROM#(.FILENAME("conv3/CONV3_36.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U35 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(35+1)-1:16*35])); 
W_ROM#(.FILENAME("conv3/CONV3_37.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U36 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(36+1)-1:16*36])); 
W_ROM#(.FILENAME("conv3/CONV3_38.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U37 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(37+1)-1:16*37])); 
W_ROM#(.FILENAME("conv3/CONV3_39.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U38 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(38+1)-1:16*38])); 
W_ROM#(.FILENAME("conv3/CONV3_40.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U39 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(39+1)-1:16*39])); 
W_ROM#(.FILENAME("conv3/CONV3_41.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U40 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(40+1)-1:16*40])); 
W_ROM#(.FILENAME("conv3/CONV3_42.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U41 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(41+1)-1:16*41])); 
W_ROM#(.FILENAME("conv3/CONV3_43.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U42 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(42+1)-1:16*42])); 
W_ROM#(.FILENAME("conv3/CONV3_44.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U43 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(43+1)-1:16*43])); 
W_ROM#(.FILENAME("conv3/CONV3_45.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U44 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(44+1)-1:16*44])); 
W_ROM#(.FILENAME("conv3/CONV3_46.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U45 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(45+1)-1:16*45])); 
W_ROM#(.FILENAME("conv3/CONV3_47.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U46 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(46+1)-1:16*46])); 
W_ROM#(.FILENAME("conv3/CONV3_48.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U47 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(47+1)-1:16*47])); 
W_ROM#(.FILENAME("conv3/CONV3_49.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U48 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(48+1)-1:16*48])); 
W_ROM#(.FILENAME("conv3/CONV3_50.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U49 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(49+1)-1:16*49])); 
W_ROM#(.FILENAME("conv3/CONV3_51.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U50 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(50+1)-1:16*50])); 
W_ROM#(.FILENAME("conv3/CONV3_52.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U51 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(51+1)-1:16*51])); 
W_ROM#(.FILENAME("conv3/CONV3_53.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U52 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(52+1)-1:16*52])); 
W_ROM#(.FILENAME("conv3/CONV3_54.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U53 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(53+1)-1:16*53])); 
W_ROM#(.FILENAME("conv3/CONV3_55.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U54 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(54+1)-1:16*54])); 
W_ROM#(.FILENAME("conv3/CONV3_56.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U55 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(55+1)-1:16*55])); 
W_ROM#(.FILENAME("conv3/CONV3_57.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U56 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(56+1)-1:16*56])); 
W_ROM#(.FILENAME("conv3/CONV3_58.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U57 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(57+1)-1:16*57])); 
W_ROM#(.FILENAME("conv3/CONV3_59.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U58 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(58+1)-1:16*58])); 
W_ROM#(.FILENAME("conv3/CONV3_60.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U59 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(59+1)-1:16*59])); 
W_ROM#(.FILENAME("conv3/CONV3_61.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U60 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(60+1)-1:16*60])); 
W_ROM#(.FILENAME("conv3/CONV3_62.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U61 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(61+1)-1:16*61])); 
W_ROM#(.FILENAME("conv3/CONV3_63.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U62 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(62+1)-1:16*62])); 
W_ROM#(.FILENAME("conv3/CONV3_64.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U63 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(63+1)-1:16*63])); 
W_ROM#(.FILENAME("conv3/CONV3_65.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U64 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(64+1)-1:16*64])); 
W_ROM#(.FILENAME("conv3/CONV3_66.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U65 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(65+1)-1:16*65])); 
W_ROM#(.FILENAME("conv3/CONV3_67.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U66 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(66+1)-1:16*66])); 
W_ROM#(.FILENAME("conv3/CONV3_68.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U67 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(67+1)-1:16*67])); 
W_ROM#(.FILENAME("conv3/CONV3_69.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U68 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(68+1)-1:16*68])); 
W_ROM#(.FILENAME("conv3/CONV3_70.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U69 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(69+1)-1:16*69])); 
W_ROM#(.FILENAME("conv3/CONV3_71.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U70 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(70+1)-1:16*70])); 
W_ROM#(.FILENAME("conv3/CONV3_72.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U71 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(71+1)-1:16*71])); 
W_ROM#(.FILENAME("conv3/CONV3_73.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U72 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(72+1)-1:16*72])); 
W_ROM#(.FILENAME("conv3/CONV3_74.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U73 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(73+1)-1:16*73])); 
W_ROM#(.FILENAME("conv3/CONV3_75.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U74 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(74+1)-1:16*74])); 
W_ROM#(.FILENAME("conv3/CONV3_76.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U75 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(75+1)-1:16*75])); 
W_ROM#(.FILENAME("conv3/CONV3_77.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U76 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(76+1)-1:16*76])); 
W_ROM#(.FILENAME("conv3/CONV3_78.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U77 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(77+1)-1:16*77])); 
W_ROM#(.FILENAME("conv3/CONV3_79.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U78 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(78+1)-1:16*78])); 
W_ROM#(.FILENAME("conv3/CONV3_80.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U79 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(79+1)-1:16*79])); 
W_ROM#(.FILENAME("conv3/CONV3_81.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U80 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(80+1)-1:16*80])); 
W_ROM#(.FILENAME("conv3/CONV3_82.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U81 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(81+1)-1:16*81])); 
W_ROM#(.FILENAME("conv3/CONV3_83.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U82 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(82+1)-1:16*82])); 
W_ROM#(.FILENAME("conv3/CONV3_84.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U83 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(83+1)-1:16*83])); 
W_ROM#(.FILENAME("conv3/CONV3_85.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U84 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(84+1)-1:16*84])); 
W_ROM#(.FILENAME("conv3/CONV3_86.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U85 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(85+1)-1:16*85])); 
W_ROM#(.FILENAME("conv3/CONV3_87.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U86 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(86+1)-1:16*86])); 
W_ROM#(.FILENAME("conv3/CONV3_88.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U87 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(87+1)-1:16*87])); 
W_ROM#(.FILENAME("conv3/CONV3_89.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U88 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(88+1)-1:16*88])); 
W_ROM#(.FILENAME("conv3/CONV3_90.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U89 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(89+1)-1:16*89])); 
W_ROM#(.FILENAME("conv3/CONV3_91.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U90 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(90+1)-1:16*90])); 
W_ROM#(.FILENAME("conv3/CONV3_92.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U91 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(91+1)-1:16*91])); 
W_ROM#(.FILENAME("conv3/CONV3_93.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U92 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(92+1)-1:16*92])); 
W_ROM#(.FILENAME("conv3/CONV3_94.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U93 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(93+1)-1:16*93])); 
W_ROM#(.FILENAME("conv3/CONV3_95.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U94 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(94+1)-1:16*94])); 
W_ROM#(.FILENAME("conv3/CONV3_96.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U95 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(95+1)-1:16*95])); 
W_ROM#(.FILENAME("conv3/CONV3_97.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U96 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(96+1)-1:16*96])); 
W_ROM#(.FILENAME("conv3/CONV3_98.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U97 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(97+1)-1:16*97])); 
W_ROM#(.FILENAME("conv3/CONV3_99.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U98 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(98+1)-1:16*98])); 
W_ROM#(.FILENAME("conv3/CONV3_100.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U99 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(99+1)-1:16*99])); 
W_ROM#(.FILENAME("conv3/CONV3_101.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U100 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(100+1)-1:16*100])); 
W_ROM#(.FILENAME("conv3/CONV3_102.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U101 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(101+1)-1:16*101])); 
W_ROM#(.FILENAME("conv3/CONV3_103.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U102 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(102+1)-1:16*102])); 
W_ROM#(.FILENAME("conv3/CONV3_104.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U103 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(103+1)-1:16*103])); 
W_ROM#(.FILENAME("conv3/CONV3_105.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U104 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(104+1)-1:16*104])); 
W_ROM#(.FILENAME("conv3/CONV3_106.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U105 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(105+1)-1:16*105])); 
W_ROM#(.FILENAME("conv3/CONV3_107.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U106 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(106+1)-1:16*106])); 
W_ROM#(.FILENAME("conv3/CONV3_108.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U107 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(107+1)-1:16*107])); 
W_ROM#(.FILENAME("conv3/CONV3_109.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U108 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(108+1)-1:16*108])); 
W_ROM#(.FILENAME("conv3/CONV3_110.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U109 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(109+1)-1:16*109])); 
W_ROM#(.FILENAME("conv3/CONV3_111.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U110 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(110+1)-1:16*110])); 
W_ROM#(.FILENAME("conv3/CONV3_112.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U111 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(111+1)-1:16*111])); 
W_ROM#(.FILENAME("conv3/CONV3_113.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U112 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(112+1)-1:16*112])); 
W_ROM#(.FILENAME("conv3/CONV3_114.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U113 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(113+1)-1:16*113])); 
W_ROM#(.FILENAME("conv3/CONV3_115.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U114 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(114+1)-1:16*114])); 
W_ROM#(.FILENAME("conv3/CONV3_116.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U115 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(115+1)-1:16*115])); 
W_ROM#(.FILENAME("conv3/CONV3_117.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U116 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(116+1)-1:16*116])); 
W_ROM#(.FILENAME("conv3/CONV3_118.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U117 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(117+1)-1:16*117])); 
W_ROM#(.FILENAME("conv3/CONV3_119.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U118 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(118+1)-1:16*118])); 
W_ROM#(.FILENAME("conv3/CONV3_120.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U119 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(119+1)-1:16*119])); 
W_ROM#(.FILENAME("conv3/CONV3_121.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U120 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(120+1)-1:16*120])); 
W_ROM#(.FILENAME("conv3/CONV3_122.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U121 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(121+1)-1:16*121])); 
W_ROM#(.FILENAME("conv3/CONV3_123.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U122 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(122+1)-1:16*122])); 
W_ROM#(.FILENAME("conv3/CONV3_124.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U123 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(123+1)-1:16*123])); 
W_ROM#(.FILENAME("conv3/CONV3_125.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U124 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(124+1)-1:16*124])); 
W_ROM#(.FILENAME("conv3/CONV3_126.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U125 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(125+1)-1:16*125])); 
W_ROM#(.FILENAME("conv3/CONV3_127.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U126 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(126+1)-1:16*126])); 
W_ROM#(.FILENAME("conv3/CONV3_128.txt"),.weight_addr_WIDTH(3),.NO_ROWS(8)) U127 (.weight_addr(weight_addr),.clk(clk),.weight_out(weight_out[16*(127+1)-1:16*127])); 


endmodule
