module conv12 #(parameter N_weight_out=256,parameter weight_addr_WIDTH=4)(weight_out_conv12,weight_addr_conv12,clk);
input wire [weight_addr_WIDTH-1:0] weight_addr_conv12;
output wire [N_weight_out*16-1:0] weight_out_conv12 ;
input clk;
W_ROM #(.FILENAME("conv12/CONV12_1.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U0 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv12/CONV12_2.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U1 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv12/CONV12_3.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U2 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv12/CONV12_4.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U3 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv12/CONV12_5.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U4 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv12/CONV12_6.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U5 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv12/CONV12_7.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U6 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv12/CONV12_8.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U7 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv12/CONV12_9.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U8 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv12/CONV12_10.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U9 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv12/CONV12_11.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U10 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv12/CONV12_12.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U11 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv12/CONV12_13.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U12 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv12/CONV12_14.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U13 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv12/CONV12_15.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U14 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv12/CONV12_16.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U15 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv12/CONV12_17.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U16 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv12/CONV12_18.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U17 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv12/CONV12_19.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U18 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv12/CONV12_20.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U19 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv12/CONV12_21.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U20 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv12/CONV12_22.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U21 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv12/CONV12_23.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U22 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv12/CONV12_24.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U23 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv12/CONV12_25.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U24 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv12/CONV12_26.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U25 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv12/CONV12_27.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U26 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv12/CONV12_28.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U27 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv12/CONV12_29.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U28 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv12/CONV12_30.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U29 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv12/CONV12_31.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U30 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv12/CONV12_32.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U31 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv12/CONV12_33.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U32 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv12/CONV12_34.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U33 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv12/CONV12_35.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U34 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv12/CONV12_36.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U35 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv12/CONV12_37.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U36 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv12/CONV12_38.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U37 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv12/CONV12_39.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U38 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv12/CONV12_40.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U39 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv12/CONV12_41.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U40 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv12/CONV12_42.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U41 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv12/CONV12_43.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U42 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv12/CONV12_44.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U43 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv12/CONV12_45.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U44 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv12/CONV12_46.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U45 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv12/CONV12_47.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U46 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv12/CONV12_48.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U47 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv12/CONV12_49.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U48 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv12/CONV12_50.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U49 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv12/CONV12_51.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U50 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv12/CONV12_52.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U51 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv12/CONV12_53.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U52 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv12/CONV12_54.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U53 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv12/CONV12_55.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U54 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv12/CONV12_56.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U55 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv12/CONV12_57.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U56 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv12/CONV12_58.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U57 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv12/CONV12_59.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U58 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv12/CONV12_60.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U59 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv12/CONV12_61.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U60 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv12/CONV12_62.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U61 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv12/CONV12_63.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U62 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv12/CONV12_64.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U63 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(63+1)-1:16*63])); 
W_ROM #(.FILENAME("conv12/CONV12_65.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U64 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(64+1)-1:16*64])); 
W_ROM #(.FILENAME("conv12/CONV12_66.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U65 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(65+1)-1:16*65])); 
W_ROM #(.FILENAME("conv12/CONV12_67.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U66 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(66+1)-1:16*66])); 
W_ROM #(.FILENAME("conv12/CONV12_68.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U67 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(67+1)-1:16*67])); 
W_ROM #(.FILENAME("conv12/CONV12_69.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U68 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(68+1)-1:16*68])); 
W_ROM #(.FILENAME("conv12/CONV12_70.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U69 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(69+1)-1:16*69])); 
W_ROM #(.FILENAME("conv12/CONV12_71.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U70 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(70+1)-1:16*70])); 
W_ROM #(.FILENAME("conv12/CONV12_72.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U71 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(71+1)-1:16*71])); 
W_ROM #(.FILENAME("conv12/CONV12_73.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U72 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(72+1)-1:16*72])); 
W_ROM #(.FILENAME("conv12/CONV12_74.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U73 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(73+1)-1:16*73])); 
W_ROM #(.FILENAME("conv12/CONV12_75.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U74 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(74+1)-1:16*74])); 
W_ROM #(.FILENAME("conv12/CONV12_76.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U75 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(75+1)-1:16*75])); 
W_ROM #(.FILENAME("conv12/CONV12_77.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U76 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(76+1)-1:16*76])); 
W_ROM #(.FILENAME("conv12/CONV12_78.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U77 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(77+1)-1:16*77])); 
W_ROM #(.FILENAME("conv12/CONV12_79.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U78 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(78+1)-1:16*78])); 
W_ROM #(.FILENAME("conv12/CONV12_80.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U79 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(79+1)-1:16*79])); 
W_ROM #(.FILENAME("conv12/CONV12_81.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U80 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(80+1)-1:16*80])); 
W_ROM #(.FILENAME("conv12/CONV12_82.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U81 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(81+1)-1:16*81])); 
W_ROM #(.FILENAME("conv12/CONV12_83.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U82 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(82+1)-1:16*82])); 
W_ROM #(.FILENAME("conv12/CONV12_84.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U83 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(83+1)-1:16*83])); 
W_ROM #(.FILENAME("conv12/CONV12_85.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U84 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(84+1)-1:16*84])); 
W_ROM #(.FILENAME("conv12/CONV12_86.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U85 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(85+1)-1:16*85])); 
W_ROM #(.FILENAME("conv12/CONV12_87.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U86 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(86+1)-1:16*86])); 
W_ROM #(.FILENAME("conv12/CONV12_88.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U87 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(87+1)-1:16*87])); 
W_ROM #(.FILENAME("conv12/CONV12_89.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U88 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(88+1)-1:16*88])); 
W_ROM #(.FILENAME("conv12/CONV12_90.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U89 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(89+1)-1:16*89])); 
W_ROM #(.FILENAME("conv12/CONV12_91.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U90 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(90+1)-1:16*90])); 
W_ROM #(.FILENAME("conv12/CONV12_92.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U91 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(91+1)-1:16*91])); 
W_ROM #(.FILENAME("conv12/CONV12_93.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U92 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(92+1)-1:16*92])); 
W_ROM #(.FILENAME("conv12/CONV12_94.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U93 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(93+1)-1:16*93])); 
W_ROM #(.FILENAME("conv12/CONV12_95.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U94 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(94+1)-1:16*94])); 
W_ROM #(.FILENAME("conv12/CONV12_96.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U95 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(95+1)-1:16*95])); 
W_ROM #(.FILENAME("conv12/CONV12_97.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U96 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(96+1)-1:16*96])); 
W_ROM #(.FILENAME("conv12/CONV12_98.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U97 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(97+1)-1:16*97])); 
W_ROM #(.FILENAME("conv12/CONV12_99.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U98 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(98+1)-1:16*98])); 
W_ROM #(.FILENAME("conv12/CONV12_100.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U99 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(99+1)-1:16*99])); 
W_ROM #(.FILENAME("conv12/CONV12_101.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U100 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(100+1)-1:16*100])); 
W_ROM #(.FILENAME("conv12/CONV12_102.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U101 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(101+1)-1:16*101])); 
W_ROM #(.FILENAME("conv12/CONV12_103.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U102 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(102+1)-1:16*102])); 
W_ROM #(.FILENAME("conv12/CONV12_104.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U103 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(103+1)-1:16*103])); 
W_ROM #(.FILENAME("conv12/CONV12_105.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U104 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(104+1)-1:16*104])); 
W_ROM #(.FILENAME("conv12/CONV12_106.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U105 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(105+1)-1:16*105])); 
W_ROM #(.FILENAME("conv12/CONV12_107.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U106 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(106+1)-1:16*106])); 
W_ROM #(.FILENAME("conv12/CONV12_108.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U107 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(107+1)-1:16*107])); 
W_ROM #(.FILENAME("conv12/CONV12_109.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U108 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(108+1)-1:16*108])); 
W_ROM #(.FILENAME("conv12/CONV12_110.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U109 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(109+1)-1:16*109])); 
W_ROM #(.FILENAME("conv12/CONV12_111.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U110 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(110+1)-1:16*110])); 
W_ROM #(.FILENAME("conv12/CONV12_112.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U111 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(111+1)-1:16*111])); 
W_ROM #(.FILENAME("conv12/CONV12_113.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U112 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(112+1)-1:16*112])); 
W_ROM #(.FILENAME("conv12/CONV12_114.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U113 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(113+1)-1:16*113])); 
W_ROM #(.FILENAME("conv12/CONV12_115.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U114 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(114+1)-1:16*114])); 
W_ROM #(.FILENAME("conv12/CONV12_116.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U115 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(115+1)-1:16*115])); 
W_ROM #(.FILENAME("conv12/CONV12_117.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U116 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(116+1)-1:16*116])); 
W_ROM #(.FILENAME("conv12/CONV12_118.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U117 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(117+1)-1:16*117])); 
W_ROM #(.FILENAME("conv12/CONV12_119.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U118 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(118+1)-1:16*118])); 
W_ROM #(.FILENAME("conv12/CONV12_120.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U119 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(119+1)-1:16*119])); 
W_ROM #(.FILENAME("conv12/CONV12_121.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U120 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(120+1)-1:16*120])); 
W_ROM #(.FILENAME("conv12/CONV12_122.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U121 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(121+1)-1:16*121])); 
W_ROM #(.FILENAME("conv12/CONV12_123.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U122 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(122+1)-1:16*122])); 
W_ROM #(.FILENAME("conv12/CONV12_124.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U123 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(123+1)-1:16*123])); 
W_ROM #(.FILENAME("conv12/CONV12_125.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U124 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(124+1)-1:16*124])); 
W_ROM #(.FILENAME("conv12/CONV12_126.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U125 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(125+1)-1:16*125])); 
W_ROM #(.FILENAME("conv12/CONV12_127.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U126 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(126+1)-1:16*126])); 
W_ROM #(.FILENAME("conv12/CONV12_128.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U127 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(127+1)-1:16*127])); 
W_ROM #(.FILENAME("conv12/CONV12_129.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U128 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(128+1)-1:16*128])); 
W_ROM #(.FILENAME("conv12/CONV12_130.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U129 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(129+1)-1:16*129])); 
W_ROM #(.FILENAME("conv12/CONV12_131.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U130 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(130+1)-1:16*130])); 
W_ROM #(.FILENAME("conv12/CONV12_132.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U131 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(131+1)-1:16*131])); 
W_ROM #(.FILENAME("conv12/CONV12_133.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U132 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(132+1)-1:16*132])); 
W_ROM #(.FILENAME("conv12/CONV12_134.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U133 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(133+1)-1:16*133])); 
W_ROM #(.FILENAME("conv12/CONV12_135.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U134 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(134+1)-1:16*134])); 
W_ROM #(.FILENAME("conv12/CONV12_136.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U135 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(135+1)-1:16*135])); 
W_ROM #(.FILENAME("conv12/CONV12_137.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U136 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(136+1)-1:16*136])); 
W_ROM #(.FILENAME("conv12/CONV12_138.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U137 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(137+1)-1:16*137])); 
W_ROM #(.FILENAME("conv12/CONV12_139.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U138 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(138+1)-1:16*138])); 
W_ROM #(.FILENAME("conv12/CONV12_140.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U139 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(139+1)-1:16*139])); 
W_ROM #(.FILENAME("conv12/CONV12_141.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U140 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(140+1)-1:16*140])); 
W_ROM #(.FILENAME("conv12/CONV12_142.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U141 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(141+1)-1:16*141])); 
W_ROM #(.FILENAME("conv12/CONV12_143.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U142 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(142+1)-1:16*142])); 
W_ROM #(.FILENAME("conv12/CONV12_144.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U143 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(143+1)-1:16*143])); 
W_ROM #(.FILENAME("conv12/CONV12_145.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U144 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(144+1)-1:16*144])); 
W_ROM #(.FILENAME("conv12/CONV12_146.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U145 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(145+1)-1:16*145])); 
W_ROM #(.FILENAME("conv12/CONV12_147.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U146 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(146+1)-1:16*146])); 
W_ROM #(.FILENAME("conv12/CONV12_148.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U147 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(147+1)-1:16*147])); 
W_ROM #(.FILENAME("conv12/CONV12_149.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U148 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(148+1)-1:16*148])); 
W_ROM #(.FILENAME("conv12/CONV12_150.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U149 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(149+1)-1:16*149])); 
W_ROM #(.FILENAME("conv12/CONV12_151.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U150 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(150+1)-1:16*150])); 
W_ROM #(.FILENAME("conv12/CONV12_152.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U151 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(151+1)-1:16*151])); 
W_ROM #(.FILENAME("conv12/CONV12_153.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U152 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(152+1)-1:16*152])); 
W_ROM #(.FILENAME("conv12/CONV12_154.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U153 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(153+1)-1:16*153])); 
W_ROM #(.FILENAME("conv12/CONV12_155.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U154 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(154+1)-1:16*154])); 
W_ROM #(.FILENAME("conv12/CONV12_156.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U155 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(155+1)-1:16*155])); 
W_ROM #(.FILENAME("conv12/CONV12_157.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U156 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(156+1)-1:16*156])); 
W_ROM #(.FILENAME("conv12/CONV12_158.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U157 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(157+1)-1:16*157])); 
W_ROM #(.FILENAME("conv12/CONV12_159.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U158 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(158+1)-1:16*158])); 
W_ROM #(.FILENAME("conv12/CONV12_160.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U159 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(159+1)-1:16*159])); 
W_ROM #(.FILENAME("conv12/CONV12_161.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U160 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(160+1)-1:16*160])); 
W_ROM #(.FILENAME("conv12/CONV12_162.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U161 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(161+1)-1:16*161])); 
W_ROM #(.FILENAME("conv12/CONV12_163.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U162 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(162+1)-1:16*162])); 
W_ROM #(.FILENAME("conv12/CONV12_164.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U163 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(163+1)-1:16*163])); 
W_ROM #(.FILENAME("conv12/CONV12_165.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U164 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(164+1)-1:16*164])); 
W_ROM #(.FILENAME("conv12/CONV12_166.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U165 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(165+1)-1:16*165])); 
W_ROM #(.FILENAME("conv12/CONV12_167.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U166 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(166+1)-1:16*166])); 
W_ROM #(.FILENAME("conv12/CONV12_168.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U167 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(167+1)-1:16*167])); 
W_ROM #(.FILENAME("conv12/CONV12_169.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U168 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(168+1)-1:16*168])); 
W_ROM #(.FILENAME("conv12/CONV12_170.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U169 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(169+1)-1:16*169])); 
W_ROM #(.FILENAME("conv12/CONV12_171.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U170 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(170+1)-1:16*170])); 
W_ROM #(.FILENAME("conv12/CONV12_172.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U171 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(171+1)-1:16*171])); 
W_ROM #(.FILENAME("conv12/CONV12_173.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U172 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(172+1)-1:16*172])); 
W_ROM #(.FILENAME("conv12/CONV12_174.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U173 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(173+1)-1:16*173])); 
W_ROM #(.FILENAME("conv12/CONV12_175.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U174 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(174+1)-1:16*174])); 
W_ROM #(.FILENAME("conv12/CONV12_176.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U175 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(175+1)-1:16*175])); 
W_ROM #(.FILENAME("conv12/CONV12_177.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U176 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(176+1)-1:16*176])); 
W_ROM #(.FILENAME("conv12/CONV12_178.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U177 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(177+1)-1:16*177])); 
W_ROM #(.FILENAME("conv12/CONV12_179.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U178 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(178+1)-1:16*178])); 
W_ROM #(.FILENAME("conv12/CONV12_180.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U179 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(179+1)-1:16*179])); 
W_ROM #(.FILENAME("conv12/CONV12_181.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U180 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(180+1)-1:16*180])); 
W_ROM #(.FILENAME("conv12/CONV12_182.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U181 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(181+1)-1:16*181])); 
W_ROM #(.FILENAME("conv12/CONV12_183.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U182 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(182+1)-1:16*182])); 
W_ROM #(.FILENAME("conv12/CONV12_184.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U183 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(183+1)-1:16*183])); 
W_ROM #(.FILENAME("conv12/CONV12_185.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U184 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(184+1)-1:16*184])); 
W_ROM #(.FILENAME("conv12/CONV12_186.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U185 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(185+1)-1:16*185])); 
W_ROM #(.FILENAME("conv12/CONV12_187.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U186 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(186+1)-1:16*186])); 
W_ROM #(.FILENAME("conv12/CONV12_188.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U187 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(187+1)-1:16*187])); 
W_ROM #(.FILENAME("conv12/CONV12_189.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U188 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(188+1)-1:16*188])); 
W_ROM #(.FILENAME("conv12/CONV12_190.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U189 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(189+1)-1:16*189])); 
W_ROM #(.FILENAME("conv12/CONV12_191.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U190 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(190+1)-1:16*190])); 
W_ROM #(.FILENAME("conv12/CONV12_192.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U191 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(191+1)-1:16*191])); 
W_ROM #(.FILENAME("conv12/CONV12_193.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U192 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(192+1)-1:16*192])); 
W_ROM #(.FILENAME("conv12/CONV12_194.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U193 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(193+1)-1:16*193])); 
W_ROM #(.FILENAME("conv12/CONV12_195.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U194 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(194+1)-1:16*194])); 
W_ROM #(.FILENAME("conv12/CONV12_196.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U195 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(195+1)-1:16*195])); 
W_ROM #(.FILENAME("conv12/CONV12_197.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U196 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(196+1)-1:16*196])); 
W_ROM #(.FILENAME("conv12/CONV12_198.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U197 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(197+1)-1:16*197])); 
W_ROM #(.FILENAME("conv12/CONV12_199.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U198 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(198+1)-1:16*198])); 
W_ROM #(.FILENAME("conv12/CONV12_200.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U199 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(199+1)-1:16*199])); 
W_ROM #(.FILENAME("conv12/CONV12_201.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U200 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(200+1)-1:16*200])); 
W_ROM #(.FILENAME("conv12/CONV12_202.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U201 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(201+1)-1:16*201])); 
W_ROM #(.FILENAME("conv12/CONV12_203.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U202 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(202+1)-1:16*202])); 
W_ROM #(.FILENAME("conv12/CONV12_204.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U203 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(203+1)-1:16*203])); 
W_ROM #(.FILENAME("conv12/CONV12_205.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U204 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(204+1)-1:16*204])); 
W_ROM #(.FILENAME("conv12/CONV12_206.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U205 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(205+1)-1:16*205])); 
W_ROM #(.FILENAME("conv12/CONV12_207.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U206 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(206+1)-1:16*206])); 
W_ROM #(.FILENAME("conv12/CONV12_208.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U207 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(207+1)-1:16*207])); 
W_ROM #(.FILENAME("conv12/CONV12_209.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U208 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(208+1)-1:16*208])); 
W_ROM #(.FILENAME("conv12/CONV12_210.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U209 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(209+1)-1:16*209])); 
W_ROM #(.FILENAME("conv12/CONV12_211.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U210 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(210+1)-1:16*210])); 
W_ROM #(.FILENAME("conv12/CONV12_212.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U211 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(211+1)-1:16*211])); 
W_ROM #(.FILENAME("conv12/CONV12_213.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U212 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(212+1)-1:16*212])); 
W_ROM #(.FILENAME("conv12/CONV12_214.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U213 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(213+1)-1:16*213])); 
W_ROM #(.FILENAME("conv12/CONV12_215.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U214 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(214+1)-1:16*214])); 
W_ROM #(.FILENAME("conv12/CONV12_216.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U215 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(215+1)-1:16*215])); 
W_ROM #(.FILENAME("conv12/CONV12_217.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U216 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(216+1)-1:16*216])); 
W_ROM #(.FILENAME("conv12/CONV12_218.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U217 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(217+1)-1:16*217])); 
W_ROM #(.FILENAME("conv12/CONV12_219.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U218 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(218+1)-1:16*218])); 
W_ROM #(.FILENAME("conv12/CONV12_220.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U219 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(219+1)-1:16*219])); 
W_ROM #(.FILENAME("conv12/CONV12_221.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U220 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(220+1)-1:16*220])); 
W_ROM #(.FILENAME("conv12/CONV12_222.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U221 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(221+1)-1:16*221])); 
W_ROM #(.FILENAME("conv12/CONV12_223.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U222 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(222+1)-1:16*222])); 
W_ROM #(.FILENAME("conv12/CONV12_224.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U223 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(223+1)-1:16*223])); 
W_ROM #(.FILENAME("conv12/CONV12_225.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U224 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(224+1)-1:16*224])); 
W_ROM #(.FILENAME("conv12/CONV12_226.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U225 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(225+1)-1:16*225])); 
W_ROM #(.FILENAME("conv12/CONV12_227.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U226 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(226+1)-1:16*226])); 
W_ROM #(.FILENAME("conv12/CONV12_228.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U227 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(227+1)-1:16*227])); 
W_ROM #(.FILENAME("conv12/CONV12_229.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U228 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(228+1)-1:16*228])); 
W_ROM #(.FILENAME("conv12/CONV12_230.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U229 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(229+1)-1:16*229])); 
W_ROM #(.FILENAME("conv12/CONV12_231.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U230 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(230+1)-1:16*230])); 
W_ROM #(.FILENAME("conv12/CONV12_232.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U231 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(231+1)-1:16*231])); 
W_ROM #(.FILENAME("conv12/CONV12_233.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U232 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(232+1)-1:16*232])); 
W_ROM #(.FILENAME("conv12/CONV12_234.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U233 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(233+1)-1:16*233])); 
W_ROM #(.FILENAME("conv12/CONV12_235.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U234 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(234+1)-1:16*234])); 
W_ROM #(.FILENAME("conv12/CONV12_236.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U235 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(235+1)-1:16*235])); 
W_ROM #(.FILENAME("conv12/CONV12_237.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U236 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(236+1)-1:16*236])); 
W_ROM #(.FILENAME("conv12/CONV12_238.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U237 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(237+1)-1:16*237])); 
W_ROM #(.FILENAME("conv12/CONV12_239.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U238 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(238+1)-1:16*238])); 
W_ROM #(.FILENAME("conv12/CONV12_240.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U239 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(239+1)-1:16*239])); 
W_ROM #(.FILENAME("conv12/CONV12_241.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U240 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(240+1)-1:16*240])); 
W_ROM #(.FILENAME("conv12/CONV12_242.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U241 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(241+1)-1:16*241])); 
W_ROM #(.FILENAME("conv12/CONV12_243.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U242 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(242+1)-1:16*242])); 
W_ROM #(.FILENAME("conv12/CONV12_244.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U243 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(243+1)-1:16*243])); 
W_ROM #(.FILENAME("conv12/CONV12_245.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U244 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(244+1)-1:16*244])); 
W_ROM #(.FILENAME("conv12/CONV12_246.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U245 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(245+1)-1:16*245])); 
W_ROM #(.FILENAME("conv12/CONV12_247.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U246 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(246+1)-1:16*246])); 
W_ROM #(.FILENAME("conv12/CONV12_248.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U247 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(247+1)-1:16*247])); 
W_ROM #(.FILENAME("conv12/CONV12_249.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U248 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(248+1)-1:16*248])); 
W_ROM #(.FILENAME("conv12/CONV12_250.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U249 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(249+1)-1:16*249])); 
W_ROM #(.FILENAME("conv12/CONV12_251.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U250 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(250+1)-1:16*250])); 
W_ROM #(.FILENAME("conv12/CONV12_252.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U251 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(251+1)-1:16*251])); 
W_ROM #(.FILENAME("conv12/CONV12_253.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U252 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(252+1)-1:16*252])); 
W_ROM #(.FILENAME("conv12/CONV12_254.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U253 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(253+1)-1:16*253])); 
W_ROM #(.FILENAME("conv12/CONV12_255.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U254 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(254+1)-1:16*254])); 
W_ROM #(.FILENAME("conv12/CONV12_256.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U255 (.weight_addr(weight_addr_conv12),.clk(clk),.weight_out(weight_out_conv12[16*(255+1)-1:16*255])); 


endmodule

