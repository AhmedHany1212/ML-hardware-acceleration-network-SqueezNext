module BIAS #(parameter value=18'b0010000000000000)(q);
output [17:0] q;

assign q=value;

endmodule
