module BIAS_layer17_60_10 #(parameter N_adder_tree=16)(q);
output wire [N_adder_tree*18-1:0] q;


BIAS #(.value(18'b000010001111100110))  U0 (.q(q[18*(0+1)-1:18*0]));
BIAS #(.value(18'b000001011010011000))  U1 (.q(q[18*(1+1)-1:18*1]));
BIAS #(.value(18'b000000101001001010))  U2 (.q(q[18*(2+1)-1:18*2]));
BIAS #(.value(18'b000001010111110110))  U3 (.q(q[18*(3+1)-1:18*3]));
BIAS #(.value(18'b000000100101100100))  U4 (.q(q[18*(4+1)-1:18*4]));
BIAS #(.value(18'b000001001101111110))  U5 (.q(q[18*(5+1)-1:18*5]));
BIAS #(.value(18'b000000011000011110))  U6 (.q(q[18*(6+1)-1:18*6]));
BIAS #(.value(18'b000001110100111110))  U7 (.q(q[18*(7+1)-1:18*7]));
BIAS #(.value(18'b000001110100011000))  U8 (.q(q[18*(8+1)-1:18*8]));
BIAS #(.value(18'b000000000010100100))  U9 (.q(q[18*(9+1)-1:18*9]));
BIAS #(.value(18'b111111001101111000))  U10 (.q(q[18*(10+1)-1:18*10]));
BIAS #(.value(18'b000000010110011100))  U11 (.q(q[18*(11+1)-1:18*11]));
BIAS #(.value(18'b000000100110011000))  U12 (.q(q[18*(12+1)-1:18*12]));
BIAS #(.value(18'b111101011010011000))  U13 (.q(q[18*(13+1)-1:18*13]));
BIAS #(.value(18'b000001000000111000))  U14 (.q(q[18*(14+1)-1:18*14]));
BIAS #(.value(18'b111111101100101100))  U15 (.q(q[18*(15+1)-1:18*15]));


endmodule
