module CONV29 #(parameter N=256,parameter weight_addr_WIDTH=5 , parameter NO_ROWS=32 )(weight_out,addr,clk);
input wire [weight_addr_WIDTH-1:0] addr;
input wire clk;
output wire [N*16-1:0] weight_out ;
W_ROM #(.FILENAME("conv29/CONV29_1.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U0 (.weight_addr(addr),.weight_out(weight_out[16*(0+1)-1:16*0]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_2.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U1 (.weight_addr(addr),.weight_out(weight_out[16*(1+1)-1:16*1]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_3.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U2 (.weight_addr(addr),.weight_out(weight_out[16*(2+1)-1:16*2]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_4.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U3 (.weight_addr(addr),.weight_out(weight_out[16*(3+1)-1:16*3]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_5.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U4 (.weight_addr(addr),.weight_out(weight_out[16*(4+1)-1:16*4]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_6.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U5 (.weight_addr(addr),.weight_out(weight_out[16*(5+1)-1:16*5]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_7.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U6 (.weight_addr(addr),.weight_out(weight_out[16*(6+1)-1:16*6]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_8.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U7 (.weight_addr(addr),.weight_out(weight_out[16*(7+1)-1:16*7]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_9.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U8 (.weight_addr(addr),.weight_out(weight_out[16*(8+1)-1:16*8]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_10.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U9 (.weight_addr(addr),.weight_out(weight_out[16*(9+1)-1:16*9]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_11.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U10 (.weight_addr(addr),.weight_out(weight_out[16*(10+1)-1:16*10]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_12.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U11 (.weight_addr(addr),.weight_out(weight_out[16*(11+1)-1:16*11]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_13.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U12 (.weight_addr(addr),.weight_out(weight_out[16*(12+1)-1:16*12]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_14.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U13 (.weight_addr(addr),.weight_out(weight_out[16*(13+1)-1:16*13]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_15.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U14 (.weight_addr(addr),.weight_out(weight_out[16*(14+1)-1:16*14]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_16.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U15 (.weight_addr(addr),.weight_out(weight_out[16*(15+1)-1:16*15]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_17.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U16 (.weight_addr(addr),.weight_out(weight_out[16*(16+1)-1:16*16]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_18.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U17 (.weight_addr(addr),.weight_out(weight_out[16*(17+1)-1:16*17]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_19.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U18 (.weight_addr(addr),.weight_out(weight_out[16*(18+1)-1:16*18]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_20.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U19 (.weight_addr(addr),.weight_out(weight_out[16*(19+1)-1:16*19]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_21.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U20 (.weight_addr(addr),.weight_out(weight_out[16*(20+1)-1:16*20]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_22.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U21 (.weight_addr(addr),.weight_out(weight_out[16*(21+1)-1:16*21]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_23.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U22 (.weight_addr(addr),.weight_out(weight_out[16*(22+1)-1:16*22]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_24.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U23 (.weight_addr(addr),.weight_out(weight_out[16*(23+1)-1:16*23]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_25.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U24 (.weight_addr(addr),.weight_out(weight_out[16*(24+1)-1:16*24]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_26.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U25 (.weight_addr(addr),.weight_out(weight_out[16*(25+1)-1:16*25]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_27.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U26 (.weight_addr(addr),.weight_out(weight_out[16*(26+1)-1:16*26]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_28.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U27 (.weight_addr(addr),.weight_out(weight_out[16*(27+1)-1:16*27]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_29.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U28 (.weight_addr(addr),.weight_out(weight_out[16*(28+1)-1:16*28]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_30.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U29 (.weight_addr(addr),.weight_out(weight_out[16*(29+1)-1:16*29]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_31.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U30 (.weight_addr(addr),.weight_out(weight_out[16*(30+1)-1:16*30]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_32.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U31 (.weight_addr(addr),.weight_out(weight_out[16*(31+1)-1:16*31]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_33.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U32 (.weight_addr(addr),.weight_out(weight_out[16*(32+1)-1:16*32]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_34.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U33 (.weight_addr(addr),.weight_out(weight_out[16*(33+1)-1:16*33]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_35.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U34 (.weight_addr(addr),.weight_out(weight_out[16*(34+1)-1:16*34]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_36.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U35 (.weight_addr(addr),.weight_out(weight_out[16*(35+1)-1:16*35]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_37.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U36 (.weight_addr(addr),.weight_out(weight_out[16*(36+1)-1:16*36]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_38.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U37 (.weight_addr(addr),.weight_out(weight_out[16*(37+1)-1:16*37]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_39.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U38 (.weight_addr(addr),.weight_out(weight_out[16*(38+1)-1:16*38]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_40.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U39 (.weight_addr(addr),.weight_out(weight_out[16*(39+1)-1:16*39]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_41.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U40 (.weight_addr(addr),.weight_out(weight_out[16*(40+1)-1:16*40]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_42.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U41 (.weight_addr(addr),.weight_out(weight_out[16*(41+1)-1:16*41]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_43.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U42 (.weight_addr(addr),.weight_out(weight_out[16*(42+1)-1:16*42]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_44.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U43 (.weight_addr(addr),.weight_out(weight_out[16*(43+1)-1:16*43]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_45.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U44 (.weight_addr(addr),.weight_out(weight_out[16*(44+1)-1:16*44]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_46.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U45 (.weight_addr(addr),.weight_out(weight_out[16*(45+1)-1:16*45]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_47.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U46 (.weight_addr(addr),.weight_out(weight_out[16*(46+1)-1:16*46]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_48.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U47 (.weight_addr(addr),.weight_out(weight_out[16*(47+1)-1:16*47]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_49.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U48 (.weight_addr(addr),.weight_out(weight_out[16*(48+1)-1:16*48]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_50.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U49 (.weight_addr(addr),.weight_out(weight_out[16*(49+1)-1:16*49]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_51.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U50 (.weight_addr(addr),.weight_out(weight_out[16*(50+1)-1:16*50]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_52.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U51 (.weight_addr(addr),.weight_out(weight_out[16*(51+1)-1:16*51]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_53.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U52 (.weight_addr(addr),.weight_out(weight_out[16*(52+1)-1:16*52]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_54.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U53 (.weight_addr(addr),.weight_out(weight_out[16*(53+1)-1:16*53]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_55.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U54 (.weight_addr(addr),.weight_out(weight_out[16*(54+1)-1:16*54]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_56.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U55 (.weight_addr(addr),.weight_out(weight_out[16*(55+1)-1:16*55]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_57.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U56 (.weight_addr(addr),.weight_out(weight_out[16*(56+1)-1:16*56]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_58.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U57 (.weight_addr(addr),.weight_out(weight_out[16*(57+1)-1:16*57]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_59.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U58 (.weight_addr(addr),.weight_out(weight_out[16*(58+1)-1:16*58]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_60.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U59 (.weight_addr(addr),.weight_out(weight_out[16*(59+1)-1:16*59]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_61.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U60 (.weight_addr(addr),.weight_out(weight_out[16*(60+1)-1:16*60]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_62.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U61 (.weight_addr(addr),.weight_out(weight_out[16*(61+1)-1:16*61]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_63.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U62 (.weight_addr(addr),.weight_out(weight_out[16*(62+1)-1:16*62]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_64.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U63 (.weight_addr(addr),.weight_out(weight_out[16*(63+1)-1:16*63]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_65.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U64 (.weight_addr(addr),.weight_out(weight_out[16*(64+1)-1:16*64]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_66.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U65 (.weight_addr(addr),.weight_out(weight_out[16*(65+1)-1:16*65]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_67.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U66 (.weight_addr(addr),.weight_out(weight_out[16*(66+1)-1:16*66]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_68.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U67 (.weight_addr(addr),.weight_out(weight_out[16*(67+1)-1:16*67]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_69.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U68 (.weight_addr(addr),.weight_out(weight_out[16*(68+1)-1:16*68]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_70.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U69 (.weight_addr(addr),.weight_out(weight_out[16*(69+1)-1:16*69]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_71.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U70 (.weight_addr(addr),.weight_out(weight_out[16*(70+1)-1:16*70]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_72.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U71 (.weight_addr(addr),.weight_out(weight_out[16*(71+1)-1:16*71]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_73.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U72 (.weight_addr(addr),.weight_out(weight_out[16*(72+1)-1:16*72]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_74.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U73 (.weight_addr(addr),.weight_out(weight_out[16*(73+1)-1:16*73]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_75.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U74 (.weight_addr(addr),.weight_out(weight_out[16*(74+1)-1:16*74]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_76.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U75 (.weight_addr(addr),.weight_out(weight_out[16*(75+1)-1:16*75]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_77.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U76 (.weight_addr(addr),.weight_out(weight_out[16*(76+1)-1:16*76]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_78.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U77 (.weight_addr(addr),.weight_out(weight_out[16*(77+1)-1:16*77]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_79.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U78 (.weight_addr(addr),.weight_out(weight_out[16*(78+1)-1:16*78]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_80.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U79 (.weight_addr(addr),.weight_out(weight_out[16*(79+1)-1:16*79]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_81.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U80 (.weight_addr(addr),.weight_out(weight_out[16*(80+1)-1:16*80]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_82.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U81 (.weight_addr(addr),.weight_out(weight_out[16*(81+1)-1:16*81]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_83.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U82 (.weight_addr(addr),.weight_out(weight_out[16*(82+1)-1:16*82]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_84.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U83 (.weight_addr(addr),.weight_out(weight_out[16*(83+1)-1:16*83]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_85.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U84 (.weight_addr(addr),.weight_out(weight_out[16*(84+1)-1:16*84]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_86.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U85 (.weight_addr(addr),.weight_out(weight_out[16*(85+1)-1:16*85]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_87.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U86 (.weight_addr(addr),.weight_out(weight_out[16*(86+1)-1:16*86]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_88.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U87 (.weight_addr(addr),.weight_out(weight_out[16*(87+1)-1:16*87]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_89.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U88 (.weight_addr(addr),.weight_out(weight_out[16*(88+1)-1:16*88]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_90.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U89 (.weight_addr(addr),.weight_out(weight_out[16*(89+1)-1:16*89]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_91.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U90 (.weight_addr(addr),.weight_out(weight_out[16*(90+1)-1:16*90]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_92.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U91 (.weight_addr(addr),.weight_out(weight_out[16*(91+1)-1:16*91]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_93.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U92 (.weight_addr(addr),.weight_out(weight_out[16*(92+1)-1:16*92]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_94.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U93 (.weight_addr(addr),.weight_out(weight_out[16*(93+1)-1:16*93]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_95.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U94 (.weight_addr(addr),.weight_out(weight_out[16*(94+1)-1:16*94]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_96.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U95 (.weight_addr(addr),.weight_out(weight_out[16*(95+1)-1:16*95]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_97.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U96 (.weight_addr(addr),.weight_out(weight_out[16*(96+1)-1:16*96]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_98.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U97 (.weight_addr(addr),.weight_out(weight_out[16*(97+1)-1:16*97]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_99.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U98 (.weight_addr(addr),.weight_out(weight_out[16*(98+1)-1:16*98]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_100.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U99 (.weight_addr(addr),.weight_out(weight_out[16*(99+1)-1:16*99]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_101.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U100 (.weight_addr(addr),.weight_out(weight_out[16*(100+1)-1:16*100]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_102.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U101 (.weight_addr(addr),.weight_out(weight_out[16*(101+1)-1:16*101]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_103.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U102 (.weight_addr(addr),.weight_out(weight_out[16*(102+1)-1:16*102]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_104.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U103 (.weight_addr(addr),.weight_out(weight_out[16*(103+1)-1:16*103]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_105.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U104 (.weight_addr(addr),.weight_out(weight_out[16*(104+1)-1:16*104]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_106.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U105 (.weight_addr(addr),.weight_out(weight_out[16*(105+1)-1:16*105]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_107.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U106 (.weight_addr(addr),.weight_out(weight_out[16*(106+1)-1:16*106]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_108.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U107 (.weight_addr(addr),.weight_out(weight_out[16*(107+1)-1:16*107]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_109.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U108 (.weight_addr(addr),.weight_out(weight_out[16*(108+1)-1:16*108]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_110.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U109 (.weight_addr(addr),.weight_out(weight_out[16*(109+1)-1:16*109]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_111.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U110 (.weight_addr(addr),.weight_out(weight_out[16*(110+1)-1:16*110]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_112.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U111 (.weight_addr(addr),.weight_out(weight_out[16*(111+1)-1:16*111]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_113.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U112 (.weight_addr(addr),.weight_out(weight_out[16*(112+1)-1:16*112]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_114.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U113 (.weight_addr(addr),.weight_out(weight_out[16*(113+1)-1:16*113]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_115.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U114 (.weight_addr(addr),.weight_out(weight_out[16*(114+1)-1:16*114]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_116.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U115 (.weight_addr(addr),.weight_out(weight_out[16*(115+1)-1:16*115]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_117.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U116 (.weight_addr(addr),.weight_out(weight_out[16*(116+1)-1:16*116]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_118.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U117 (.weight_addr(addr),.weight_out(weight_out[16*(117+1)-1:16*117]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_119.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U118 (.weight_addr(addr),.weight_out(weight_out[16*(118+1)-1:16*118]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_120.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U119 (.weight_addr(addr),.weight_out(weight_out[16*(119+1)-1:16*119]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_121.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U120 (.weight_addr(addr),.weight_out(weight_out[16*(120+1)-1:16*120]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_122.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U121 (.weight_addr(addr),.weight_out(weight_out[16*(121+1)-1:16*121]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_123.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U122 (.weight_addr(addr),.weight_out(weight_out[16*(122+1)-1:16*122]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_124.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U123 (.weight_addr(addr),.weight_out(weight_out[16*(123+1)-1:16*123]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_125.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U124 (.weight_addr(addr),.weight_out(weight_out[16*(124+1)-1:16*124]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_126.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U125 (.weight_addr(addr),.weight_out(weight_out[16*(125+1)-1:16*125]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_127.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U126 (.weight_addr(addr),.weight_out(weight_out[16*(126+1)-1:16*126]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_128.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U127 (.weight_addr(addr),.weight_out(weight_out[16*(127+1)-1:16*127]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_129.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U128 (.weight_addr(addr),.weight_out(weight_out[16*(128+1)-1:16*128]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_130.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U129 (.weight_addr(addr),.weight_out(weight_out[16*(129+1)-1:16*129]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_131.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U130 (.weight_addr(addr),.weight_out(weight_out[16*(130+1)-1:16*130]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_132.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U131 (.weight_addr(addr),.weight_out(weight_out[16*(131+1)-1:16*131]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_133.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U132 (.weight_addr(addr),.weight_out(weight_out[16*(132+1)-1:16*132]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_134.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U133 (.weight_addr(addr),.weight_out(weight_out[16*(133+1)-1:16*133]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_135.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U134 (.weight_addr(addr),.weight_out(weight_out[16*(134+1)-1:16*134]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_136.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U135 (.weight_addr(addr),.weight_out(weight_out[16*(135+1)-1:16*135]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_137.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U136 (.weight_addr(addr),.weight_out(weight_out[16*(136+1)-1:16*136]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_138.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U137 (.weight_addr(addr),.weight_out(weight_out[16*(137+1)-1:16*137]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_139.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U138 (.weight_addr(addr),.weight_out(weight_out[16*(138+1)-1:16*138]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_140.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U139 (.weight_addr(addr),.weight_out(weight_out[16*(139+1)-1:16*139]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_141.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U140 (.weight_addr(addr),.weight_out(weight_out[16*(140+1)-1:16*140]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_142.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U141 (.weight_addr(addr),.weight_out(weight_out[16*(141+1)-1:16*141]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_143.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U142 (.weight_addr(addr),.weight_out(weight_out[16*(142+1)-1:16*142]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_144.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U143 (.weight_addr(addr),.weight_out(weight_out[16*(143+1)-1:16*143]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_145.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U144 (.weight_addr(addr),.weight_out(weight_out[16*(144+1)-1:16*144]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_146.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U145 (.weight_addr(addr),.weight_out(weight_out[16*(145+1)-1:16*145]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_147.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U146 (.weight_addr(addr),.weight_out(weight_out[16*(146+1)-1:16*146]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_148.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U147 (.weight_addr(addr),.weight_out(weight_out[16*(147+1)-1:16*147]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_149.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U148 (.weight_addr(addr),.weight_out(weight_out[16*(148+1)-1:16*148]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_150.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U149 (.weight_addr(addr),.weight_out(weight_out[16*(149+1)-1:16*149]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_151.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U150 (.weight_addr(addr),.weight_out(weight_out[16*(150+1)-1:16*150]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_152.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U151 (.weight_addr(addr),.weight_out(weight_out[16*(151+1)-1:16*151]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_153.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U152 (.weight_addr(addr),.weight_out(weight_out[16*(152+1)-1:16*152]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_154.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U153 (.weight_addr(addr),.weight_out(weight_out[16*(153+1)-1:16*153]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_155.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U154 (.weight_addr(addr),.weight_out(weight_out[16*(154+1)-1:16*154]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_156.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U155 (.weight_addr(addr),.weight_out(weight_out[16*(155+1)-1:16*155]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_157.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U156 (.weight_addr(addr),.weight_out(weight_out[16*(156+1)-1:16*156]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_158.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U157 (.weight_addr(addr),.weight_out(weight_out[16*(157+1)-1:16*157]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_159.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U158 (.weight_addr(addr),.weight_out(weight_out[16*(158+1)-1:16*158]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_160.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U159 (.weight_addr(addr),.weight_out(weight_out[16*(159+1)-1:16*159]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_161.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U160 (.weight_addr(addr),.weight_out(weight_out[16*(160+1)-1:16*160]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_162.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U161 (.weight_addr(addr),.weight_out(weight_out[16*(161+1)-1:16*161]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_163.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U162 (.weight_addr(addr),.weight_out(weight_out[16*(162+1)-1:16*162]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_164.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U163 (.weight_addr(addr),.weight_out(weight_out[16*(163+1)-1:16*163]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_165.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U164 (.weight_addr(addr),.weight_out(weight_out[16*(164+1)-1:16*164]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_166.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U165 (.weight_addr(addr),.weight_out(weight_out[16*(165+1)-1:16*165]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_167.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U166 (.weight_addr(addr),.weight_out(weight_out[16*(166+1)-1:16*166]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_168.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U167 (.weight_addr(addr),.weight_out(weight_out[16*(167+1)-1:16*167]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_169.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U168 (.weight_addr(addr),.weight_out(weight_out[16*(168+1)-1:16*168]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_170.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U169 (.weight_addr(addr),.weight_out(weight_out[16*(169+1)-1:16*169]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_171.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U170 (.weight_addr(addr),.weight_out(weight_out[16*(170+1)-1:16*170]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_172.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U171 (.weight_addr(addr),.weight_out(weight_out[16*(171+1)-1:16*171]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_173.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U172 (.weight_addr(addr),.weight_out(weight_out[16*(172+1)-1:16*172]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_174.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U173 (.weight_addr(addr),.weight_out(weight_out[16*(173+1)-1:16*173]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_175.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U174 (.weight_addr(addr),.weight_out(weight_out[16*(174+1)-1:16*174]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_176.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U175 (.weight_addr(addr),.weight_out(weight_out[16*(175+1)-1:16*175]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_177.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U176 (.weight_addr(addr),.weight_out(weight_out[16*(176+1)-1:16*176]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_178.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U177 (.weight_addr(addr),.weight_out(weight_out[16*(177+1)-1:16*177]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_179.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U178 (.weight_addr(addr),.weight_out(weight_out[16*(178+1)-1:16*178]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_180.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U179 (.weight_addr(addr),.weight_out(weight_out[16*(179+1)-1:16*179]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_181.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U180 (.weight_addr(addr),.weight_out(weight_out[16*(180+1)-1:16*180]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_182.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U181 (.weight_addr(addr),.weight_out(weight_out[16*(181+1)-1:16*181]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_183.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U182 (.weight_addr(addr),.weight_out(weight_out[16*(182+1)-1:16*182]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_184.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U183 (.weight_addr(addr),.weight_out(weight_out[16*(183+1)-1:16*183]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_185.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U184 (.weight_addr(addr),.weight_out(weight_out[16*(184+1)-1:16*184]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_186.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U185 (.weight_addr(addr),.weight_out(weight_out[16*(185+1)-1:16*185]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_187.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U186 (.weight_addr(addr),.weight_out(weight_out[16*(186+1)-1:16*186]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_188.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U187 (.weight_addr(addr),.weight_out(weight_out[16*(187+1)-1:16*187]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_189.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U188 (.weight_addr(addr),.weight_out(weight_out[16*(188+1)-1:16*188]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_190.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U189 (.weight_addr(addr),.weight_out(weight_out[16*(189+1)-1:16*189]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_191.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U190 (.weight_addr(addr),.weight_out(weight_out[16*(190+1)-1:16*190]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_192.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U191 (.weight_addr(addr),.weight_out(weight_out[16*(191+1)-1:16*191]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_193.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U192 (.weight_addr(addr),.weight_out(weight_out[16*(192+1)-1:16*192]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_194.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U193 (.weight_addr(addr),.weight_out(weight_out[16*(193+1)-1:16*193]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_195.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U194 (.weight_addr(addr),.weight_out(weight_out[16*(194+1)-1:16*194]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_196.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U195 (.weight_addr(addr),.weight_out(weight_out[16*(195+1)-1:16*195]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_197.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U196 (.weight_addr(addr),.weight_out(weight_out[16*(196+1)-1:16*196]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_198.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U197 (.weight_addr(addr),.weight_out(weight_out[16*(197+1)-1:16*197]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_199.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U198 (.weight_addr(addr),.weight_out(weight_out[16*(198+1)-1:16*198]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_200.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U199 (.weight_addr(addr),.weight_out(weight_out[16*(199+1)-1:16*199]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_201.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U200 (.weight_addr(addr),.weight_out(weight_out[16*(200+1)-1:16*200]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_202.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U201 (.weight_addr(addr),.weight_out(weight_out[16*(201+1)-1:16*201]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_203.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U202 (.weight_addr(addr),.weight_out(weight_out[16*(202+1)-1:16*202]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_204.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U203 (.weight_addr(addr),.weight_out(weight_out[16*(203+1)-1:16*203]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_205.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U204 (.weight_addr(addr),.weight_out(weight_out[16*(204+1)-1:16*204]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_206.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U205 (.weight_addr(addr),.weight_out(weight_out[16*(205+1)-1:16*205]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_207.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U206 (.weight_addr(addr),.weight_out(weight_out[16*(206+1)-1:16*206]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_208.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U207 (.weight_addr(addr),.weight_out(weight_out[16*(207+1)-1:16*207]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_209.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U208 (.weight_addr(addr),.weight_out(weight_out[16*(208+1)-1:16*208]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_210.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U209 (.weight_addr(addr),.weight_out(weight_out[16*(209+1)-1:16*209]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_211.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U210 (.weight_addr(addr),.weight_out(weight_out[16*(210+1)-1:16*210]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_212.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U211 (.weight_addr(addr),.weight_out(weight_out[16*(211+1)-1:16*211]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_213.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U212 (.weight_addr(addr),.weight_out(weight_out[16*(212+1)-1:16*212]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_214.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U213 (.weight_addr(addr),.weight_out(weight_out[16*(213+1)-1:16*213]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_215.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U214 (.weight_addr(addr),.weight_out(weight_out[16*(214+1)-1:16*214]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_216.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U215 (.weight_addr(addr),.weight_out(weight_out[16*(215+1)-1:16*215]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_217.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U216 (.weight_addr(addr),.weight_out(weight_out[16*(216+1)-1:16*216]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_218.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U217 (.weight_addr(addr),.weight_out(weight_out[16*(217+1)-1:16*217]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_219.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U218 (.weight_addr(addr),.weight_out(weight_out[16*(218+1)-1:16*218]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_220.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U219 (.weight_addr(addr),.weight_out(weight_out[16*(219+1)-1:16*219]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_221.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U220 (.weight_addr(addr),.weight_out(weight_out[16*(220+1)-1:16*220]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_222.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U221 (.weight_addr(addr),.weight_out(weight_out[16*(221+1)-1:16*221]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_223.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U222 (.weight_addr(addr),.weight_out(weight_out[16*(222+1)-1:16*222]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_224.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U223 (.weight_addr(addr),.weight_out(weight_out[16*(223+1)-1:16*223]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_225.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U224 (.weight_addr(addr),.weight_out(weight_out[16*(224+1)-1:16*224]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_226.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U225 (.weight_addr(addr),.weight_out(weight_out[16*(225+1)-1:16*225]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_227.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U226 (.weight_addr(addr),.weight_out(weight_out[16*(226+1)-1:16*226]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_228.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U227 (.weight_addr(addr),.weight_out(weight_out[16*(227+1)-1:16*227]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_229.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U228 (.weight_addr(addr),.weight_out(weight_out[16*(228+1)-1:16*228]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_230.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U229 (.weight_addr(addr),.weight_out(weight_out[16*(229+1)-1:16*229]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_231.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U230 (.weight_addr(addr),.weight_out(weight_out[16*(230+1)-1:16*230]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_232.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U231 (.weight_addr(addr),.weight_out(weight_out[16*(231+1)-1:16*231]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_233.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U232 (.weight_addr(addr),.weight_out(weight_out[16*(232+1)-1:16*232]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_234.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U233 (.weight_addr(addr),.weight_out(weight_out[16*(233+1)-1:16*233]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_235.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U234 (.weight_addr(addr),.weight_out(weight_out[16*(234+1)-1:16*234]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_236.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U235 (.weight_addr(addr),.weight_out(weight_out[16*(235+1)-1:16*235]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_237.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U236 (.weight_addr(addr),.weight_out(weight_out[16*(236+1)-1:16*236]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_238.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U237 (.weight_addr(addr),.weight_out(weight_out[16*(237+1)-1:16*237]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_239.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U238 (.weight_addr(addr),.weight_out(weight_out[16*(238+1)-1:16*238]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_240.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U239 (.weight_addr(addr),.weight_out(weight_out[16*(239+1)-1:16*239]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_241.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U240 (.weight_addr(addr),.weight_out(weight_out[16*(240+1)-1:16*240]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_242.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U241 (.weight_addr(addr),.weight_out(weight_out[16*(241+1)-1:16*241]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_243.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U242 (.weight_addr(addr),.weight_out(weight_out[16*(242+1)-1:16*242]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_244.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U243 (.weight_addr(addr),.weight_out(weight_out[16*(243+1)-1:16*243]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_245.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U244 (.weight_addr(addr),.weight_out(weight_out[16*(244+1)-1:16*244]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_246.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U245 (.weight_addr(addr),.weight_out(weight_out[16*(245+1)-1:16*245]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_247.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U246 (.weight_addr(addr),.weight_out(weight_out[16*(246+1)-1:16*246]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_248.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U247 (.weight_addr(addr),.weight_out(weight_out[16*(247+1)-1:16*247]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_249.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U248 (.weight_addr(addr),.weight_out(weight_out[16*(248+1)-1:16*248]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_250.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U249 (.weight_addr(addr),.weight_out(weight_out[16*(249+1)-1:16*249]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_251.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U250 (.weight_addr(addr),.weight_out(weight_out[16*(250+1)-1:16*250]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_252.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U251 (.weight_addr(addr),.weight_out(weight_out[16*(251+1)-1:16*251]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_253.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U252 (.weight_addr(addr),.weight_out(weight_out[16*(252+1)-1:16*252]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_254.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U253 (.weight_addr(addr),.weight_out(weight_out[16*(253+1)-1:16*253]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_255.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U254 (.weight_addr(addr),.weight_out(weight_out[16*(254+1)-1:16*254]),.clk(clk)); 
W_ROM #(.FILENAME("conv29/CONV29_256.txt"),.weight_addr_WIDTH(weight_addr_WIDTH),.NO_ROWS(NO_ROWS)) U255 (.weight_addr(addr),.weight_out(weight_out[16*(255+1)-1:16*255]),.clk(clk)); 
endmodule
