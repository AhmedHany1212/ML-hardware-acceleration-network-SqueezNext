module BIAS_layer17_65_1 #(parameter N_adder_tree=16)(q);
output wire [N_adder_tree*18-1:0] q;


BIAS #(.value(18'b111111110110000000))  U0 (.q(q[18*(0+1)-1:18*0]));
BIAS #(.value(18'b000000001010001000))  U1 (.q(q[18*(1+1)-1:18*1]));
BIAS #(.value(18'b000000011111111110))  U2 (.q(q[18*(2+1)-1:18*2]));
BIAS #(.value(18'b111111011010110010))  U3 (.q(q[18*(3+1)-1:18*3]));
BIAS #(.value(18'b111111011001111100))  U4 (.q(q[18*(4+1)-1:18*4]));
BIAS #(.value(18'b000000101000000010))  U5 (.q(q[18*(5+1)-1:18*5]));
BIAS #(.value(18'b111111101101111110))  U6 (.q(q[18*(6+1)-1:18*6]));
BIAS #(.value(18'b111111101010010110))  U7 (.q(q[18*(7+1)-1:18*7]));
BIAS #(.value(18'b000000100000011110))  U8 (.q(q[18*(8+1)-1:18*8]));
BIAS #(.value(18'b111111111000011100))  U9 (.q(q[18*(9+1)-1:18*9]));
BIAS #(.value(18'b000000001011110110))  U10 (.q(q[18*(10+1)-1:18*10]));
BIAS #(.value(18'b000000100100100010))  U11 (.q(q[18*(11+1)-1:18*11]));
BIAS #(.value(18'b000000010101110110))  U12 (.q(q[18*(12+1)-1:18*12]));
BIAS #(.value(18'b000000101000111110))  U13 (.q(q[18*(13+1)-1:18*13]));
BIAS #(.value(18'b000000011011000100))  U14 (.q(q[18*(14+1)-1:18*14]));
BIAS #(.value(18'b111111010110011100))  U15 (.q(q[18*(15+1)-1:18*15]));


endmodule
