module CONV6 #(parameter N=64,parameter ADDR_WIDTH=4)(addr,clk,q);
input wire [ADDR_WIDTH-1:0] addr;
output wire [N*16-1:0] q ;
input clk;

W_ROM #(.FILENAME("conv6/CONV6_1.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U0 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv6/CONV6_2.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U1 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv6/CONV6_3.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U2 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv6/CONV6_4.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U3 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv6/CONV6_5.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U4 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv6/CONV6_6.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U5 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv6/CONV6_7.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U6 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv6/CONV6_8.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U7 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv6/CONV6_9.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U8 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv6/CONV6_10.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U9 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv6/CONV6_11.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U10 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv6/CONV6_12.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U11 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv6/CONV6_13.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U12 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv6/CONV6_14.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U13 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv6/CONV6_15.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U14 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv6/CONV6_16.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U15 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv6/CONV6_17.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U16 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv6/CONV6_18.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U17 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv6/CONV6_19.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U18 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv6/CONV6_20.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U19 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv6/CONV6_21.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U20 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv6/CONV6_22.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U21 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv6/CONV6_23.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U22 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv6/CONV6_24.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U23 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv6/CONV6_25.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U24 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv6/CONV6_26.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U25 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv6/CONV6_27.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U26 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv6/CONV6_28.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U27 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv6/CONV6_29.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U28 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv6/CONV6_30.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U29 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv6/CONV6_31.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U30 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv6/CONV6_32.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U31 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv6/CONV6_33.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U32 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv6/CONV6_34.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U33 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv6/CONV6_35.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U34 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv6/CONV6_36.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U35 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv6/CONV6_37.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U36 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv6/CONV6_38.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U37 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv6/CONV6_39.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U38 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv6/CONV6_40.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U39 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv6/CONV6_41.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U40 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv6/CONV6_42.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U41 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv6/CONV6_43.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U42 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv6/CONV6_44.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U43 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv6/CONV6_45.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U44 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv6/CONV6_46.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U45 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv6/CONV6_47.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U46 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv6/CONV6_48.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U47 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv6/CONV6_49.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U48 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv6/CONV6_50.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U49 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv6/CONV6_51.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U50 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv6/CONV6_52.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U51 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv6/CONV6_53.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U52 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv6/CONV6_54.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U53 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv6/CONV6_55.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U54 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv6/CONV6_56.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U55 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv6/CONV6_57.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U56 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv6/CONV6_58.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U57 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv6/CONV6_59.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U58 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv6/CONV6_60.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U59 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv6/CONV6_61.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U60 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv6/CONV6_62.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U61 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv6/CONV6_63.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U62 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv6/CONV6_64.txt"),.weight_addr_WIDTH(4),.NO_ROWS(14)) U63 (.weight_addr(addr),.clk(clk),.weight_out(q[16*(63+1)-1:16*63])); 



endmodule
