module conv11 #(parameter N_weight_out=256,parameter weight_addr_WIDTH=3)(weight_out_conv11,weight_addr_conv11,clk);
input wire [weight_addr_WIDTH-1:0] weight_addr_conv11;
output wire [N_weight_out*16-1:0] weight_out_conv11 ;
input clk;
W_ROM #(.FILENAME("conv11/CONV11_1.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U0 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(0+1)-1:16*0])); 
W_ROM #(.FILENAME("conv11/CONV11_2.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U1 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(1+1)-1:16*1])); 
W_ROM #(.FILENAME("conv11/CONV11_3.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U2 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(2+1)-1:16*2])); 
W_ROM #(.FILENAME("conv11/CONV11_4.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U3 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(3+1)-1:16*3])); 
W_ROM #(.FILENAME("conv11/CONV11_5.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U4 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(4+1)-1:16*4])); 
W_ROM #(.FILENAME("conv11/CONV11_6.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U5 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(5+1)-1:16*5])); 
W_ROM #(.FILENAME("conv11/CONV11_7.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U6 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(6+1)-1:16*6])); 
W_ROM #(.FILENAME("conv11/CONV11_8.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U7 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(7+1)-1:16*7])); 
W_ROM #(.FILENAME("conv11/CONV11_9.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U8 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(8+1)-1:16*8])); 
W_ROM #(.FILENAME("conv11/CONV11_10.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U9 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(9+1)-1:16*9])); 
W_ROM #(.FILENAME("conv11/CONV11_11.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U10 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(10+1)-1:16*10])); 
W_ROM #(.FILENAME("conv11/CONV11_12.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U11 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(11+1)-1:16*11])); 
W_ROM #(.FILENAME("conv11/CONV11_13.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U12 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(12+1)-1:16*12])); 
W_ROM #(.FILENAME("conv11/CONV11_14.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U13 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(13+1)-1:16*13])); 
W_ROM #(.FILENAME("conv11/CONV11_15.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U14 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(14+1)-1:16*14])); 
W_ROM #(.FILENAME("conv11/CONV11_16.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U15 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(15+1)-1:16*15])); 
W_ROM #(.FILENAME("conv11/CONV11_17.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U16 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(16+1)-1:16*16])); 
W_ROM #(.FILENAME("conv11/CONV11_18.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U17 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(17+1)-1:16*17])); 
W_ROM #(.FILENAME("conv11/CONV11_19.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U18 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(18+1)-1:16*18])); 
W_ROM #(.FILENAME("conv11/CONV11_20.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U19 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(19+1)-1:16*19])); 
W_ROM #(.FILENAME("conv11/CONV11_21.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U20 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(20+1)-1:16*20])); 
W_ROM #(.FILENAME("conv11/CONV11_22.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U21 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(21+1)-1:16*21])); 
W_ROM #(.FILENAME("conv11/CONV11_23.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U22 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(22+1)-1:16*22])); 
W_ROM #(.FILENAME("conv11/CONV11_24.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U23 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(23+1)-1:16*23])); 
W_ROM #(.FILENAME("conv11/CONV11_25.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U24 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(24+1)-1:16*24])); 
W_ROM #(.FILENAME("conv11/CONV11_26.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U25 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(25+1)-1:16*25])); 
W_ROM #(.FILENAME("conv11/CONV11_27.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U26 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(26+1)-1:16*26])); 
W_ROM #(.FILENAME("conv11/CONV11_28.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U27 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(27+1)-1:16*27])); 
W_ROM #(.FILENAME("conv11/CONV11_29.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U28 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(28+1)-1:16*28])); 
W_ROM #(.FILENAME("conv11/CONV11_30.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U29 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(29+1)-1:16*29])); 
W_ROM #(.FILENAME("conv11/CONV11_31.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U30 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(30+1)-1:16*30])); 
W_ROM #(.FILENAME("conv11/CONV11_32.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U31 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(31+1)-1:16*31])); 
W_ROM #(.FILENAME("conv11/CONV11_33.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U32 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(32+1)-1:16*32])); 
W_ROM #(.FILENAME("conv11/CONV11_34.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U33 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(33+1)-1:16*33])); 
W_ROM #(.FILENAME("conv11/CONV11_35.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U34 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(34+1)-1:16*34])); 
W_ROM #(.FILENAME("conv11/CONV11_36.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U35 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(35+1)-1:16*35])); 
W_ROM #(.FILENAME("conv11/CONV11_37.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U36 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(36+1)-1:16*36])); 
W_ROM #(.FILENAME("conv11/CONV11_38.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U37 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(37+1)-1:16*37])); 
W_ROM #(.FILENAME("conv11/CONV11_39.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U38 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(38+1)-1:16*38])); 
W_ROM #(.FILENAME("conv11/CONV11_40.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U39 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(39+1)-1:16*39])); 
W_ROM #(.FILENAME("conv11/CONV11_41.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U40 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(40+1)-1:16*40])); 
W_ROM #(.FILENAME("conv11/CONV11_42.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U41 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(41+1)-1:16*41])); 
W_ROM #(.FILENAME("conv11/CONV11_43.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U42 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(42+1)-1:16*42])); 
W_ROM #(.FILENAME("conv11/CONV11_44.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U43 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(43+1)-1:16*43])); 
W_ROM #(.FILENAME("conv11/CONV11_45.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U44 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(44+1)-1:16*44])); 
W_ROM #(.FILENAME("conv11/CONV11_46.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U45 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(45+1)-1:16*45])); 
W_ROM #(.FILENAME("conv11/CONV11_47.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U46 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(46+1)-1:16*46])); 
W_ROM #(.FILENAME("conv11/CONV11_48.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U47 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(47+1)-1:16*47])); 
W_ROM #(.FILENAME("conv11/CONV11_49.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U48 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(48+1)-1:16*48])); 
W_ROM #(.FILENAME("conv11/CONV11_50.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U49 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(49+1)-1:16*49])); 
W_ROM #(.FILENAME("conv11/CONV11_51.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U50 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(50+1)-1:16*50])); 
W_ROM #(.FILENAME("conv11/CONV11_52.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U51 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(51+1)-1:16*51])); 
W_ROM #(.FILENAME("conv11/CONV11_53.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U52 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(52+1)-1:16*52])); 
W_ROM #(.FILENAME("conv11/CONV11_54.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U53 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(53+1)-1:16*53])); 
W_ROM #(.FILENAME("conv11/CONV11_55.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U54 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(54+1)-1:16*54])); 
W_ROM #(.FILENAME("conv11/CONV11_56.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U55 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(55+1)-1:16*55])); 
W_ROM #(.FILENAME("conv11/CONV11_57.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U56 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(56+1)-1:16*56])); 
W_ROM #(.FILENAME("conv11/CONV11_58.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U57 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(57+1)-1:16*57])); 
W_ROM #(.FILENAME("conv11/CONV11_59.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U58 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(58+1)-1:16*58])); 
W_ROM #(.FILENAME("conv11/CONV11_60.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U59 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(59+1)-1:16*59])); 
W_ROM #(.FILENAME("conv11/CONV11_61.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U60 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(60+1)-1:16*60])); 
W_ROM #(.FILENAME("conv11/CONV11_62.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U61 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(61+1)-1:16*61])); 
W_ROM #(.FILENAME("conv11/CONV11_63.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U62 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(62+1)-1:16*62])); 
W_ROM #(.FILENAME("conv11/CONV11_64.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U63 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(63+1)-1:16*63])); 
W_ROM #(.FILENAME("conv11/CONV11_65.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U64 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(64+1)-1:16*64])); 
W_ROM #(.FILENAME("conv11/CONV11_66.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U65 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(65+1)-1:16*65])); 
W_ROM #(.FILENAME("conv11/CONV11_67.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U66 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(66+1)-1:16*66])); 
W_ROM #(.FILENAME("conv11/CONV11_68.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U67 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(67+1)-1:16*67])); 
W_ROM #(.FILENAME("conv11/CONV11_69.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U68 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(68+1)-1:16*68])); 
W_ROM #(.FILENAME("conv11/CONV11_70.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U69 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(69+1)-1:16*69])); 
W_ROM #(.FILENAME("conv11/CONV11_71.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U70 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(70+1)-1:16*70])); 
W_ROM #(.FILENAME("conv11/CONV11_72.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U71 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(71+1)-1:16*71])); 
W_ROM #(.FILENAME("conv11/CONV11_73.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U72 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(72+1)-1:16*72])); 
W_ROM #(.FILENAME("conv11/CONV11_74.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U73 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(73+1)-1:16*73])); 
W_ROM #(.FILENAME("conv11/CONV11_75.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U74 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(74+1)-1:16*74])); 
W_ROM #(.FILENAME("conv11/CONV11_76.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U75 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(75+1)-1:16*75])); 
W_ROM #(.FILENAME("conv11/CONV11_77.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U76 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(76+1)-1:16*76])); 
W_ROM #(.FILENAME("conv11/CONV11_78.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U77 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(77+1)-1:16*77])); 
W_ROM #(.FILENAME("conv11/CONV11_79.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U78 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(78+1)-1:16*78])); 
W_ROM #(.FILENAME("conv11/CONV11_80.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U79 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(79+1)-1:16*79])); 
W_ROM #(.FILENAME("conv11/CONV11_81.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U80 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(80+1)-1:16*80])); 
W_ROM #(.FILENAME("conv11/CONV11_82.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U81 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(81+1)-1:16*81])); 
W_ROM #(.FILENAME("conv11/CONV11_83.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U82 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(82+1)-1:16*82])); 
W_ROM #(.FILENAME("conv11/CONV11_84.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U83 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(83+1)-1:16*83])); 
W_ROM #(.FILENAME("conv11/CONV11_85.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U84 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(84+1)-1:16*84])); 
W_ROM #(.FILENAME("conv11/CONV11_86.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U85 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(85+1)-1:16*85])); 
W_ROM #(.FILENAME("conv11/CONV11_87.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U86 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(86+1)-1:16*86])); 
W_ROM #(.FILENAME("conv11/CONV11_88.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U87 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(87+1)-1:16*87])); 
W_ROM #(.FILENAME("conv11/CONV11_89.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U88 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(88+1)-1:16*88])); 
W_ROM #(.FILENAME("conv11/CONV11_90.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U89 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(89+1)-1:16*89])); 
W_ROM #(.FILENAME("conv11/CONV11_91.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U90 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(90+1)-1:16*90])); 
W_ROM #(.FILENAME("conv11/CONV11_92.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U91 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(91+1)-1:16*91])); 
W_ROM #(.FILENAME("conv11/CONV11_93.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U92 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(92+1)-1:16*92])); 
W_ROM #(.FILENAME("conv11/CONV11_94.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U93 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(93+1)-1:16*93])); 
W_ROM #(.FILENAME("conv11/CONV11_95.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U94 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(94+1)-1:16*94])); 
W_ROM #(.FILENAME("conv11/CONV11_96.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U95 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(95+1)-1:16*95])); 
W_ROM #(.FILENAME("conv11/CONV11_97.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U96 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(96+1)-1:16*96])); 
W_ROM #(.FILENAME("conv11/CONV11_98.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U97 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(97+1)-1:16*97])); 
W_ROM #(.FILENAME("conv11/CONV11_99.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U98 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(98+1)-1:16*98])); 
W_ROM #(.FILENAME("conv11/CONV11_100.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U99 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(99+1)-1:16*99])); 
W_ROM #(.FILENAME("conv11/CONV11_101.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U100 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(100+1)-1:16*100])); 
W_ROM #(.FILENAME("conv11/CONV11_102.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U101 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(101+1)-1:16*101])); 
W_ROM #(.FILENAME("conv11/CONV11_103.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U102 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(102+1)-1:16*102])); 
W_ROM #(.FILENAME("conv11/CONV11_104.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U103 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(103+1)-1:16*103])); 
W_ROM #(.FILENAME("conv11/CONV11_105.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U104 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(104+1)-1:16*104])); 
W_ROM #(.FILENAME("conv11/CONV11_106.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U105 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(105+1)-1:16*105])); 
W_ROM #(.FILENAME("conv11/CONV11_107.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U106 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(106+1)-1:16*106])); 
W_ROM #(.FILENAME("conv11/CONV11_108.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U107 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(107+1)-1:16*107])); 
W_ROM #(.FILENAME("conv11/CONV11_109.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U108 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(108+1)-1:16*108])); 
W_ROM #(.FILENAME("conv11/CONV11_110.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U109 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(109+1)-1:16*109])); 
W_ROM #(.FILENAME("conv11/CONV11_111.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U110 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(110+1)-1:16*110])); 
W_ROM #(.FILENAME("conv11/CONV11_112.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U111 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(111+1)-1:16*111])); 
W_ROM #(.FILENAME("conv11/CONV11_113.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U112 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(112+1)-1:16*112])); 
W_ROM #(.FILENAME("conv11/CONV11_114.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U113 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(113+1)-1:16*113])); 
W_ROM #(.FILENAME("conv11/CONV11_115.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U114 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(114+1)-1:16*114])); 
W_ROM #(.FILENAME("conv11/CONV11_116.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U115 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(115+1)-1:16*115])); 
W_ROM #(.FILENAME("conv11/CONV11_117.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U116 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(116+1)-1:16*116])); 
W_ROM #(.FILENAME("conv11/CONV11_118.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U117 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(117+1)-1:16*117])); 
W_ROM #(.FILENAME("conv11/CONV11_119.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U118 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(118+1)-1:16*118])); 
W_ROM #(.FILENAME("conv11/CONV11_120.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U119 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(119+1)-1:16*119])); 
W_ROM #(.FILENAME("conv11/CONV11_121.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U120 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(120+1)-1:16*120])); 
W_ROM #(.FILENAME("conv11/CONV11_122.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U121 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(121+1)-1:16*121])); 
W_ROM #(.FILENAME("conv11/CONV11_123.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U122 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(122+1)-1:16*122])); 
W_ROM #(.FILENAME("conv11/CONV11_124.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U123 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(123+1)-1:16*123])); 
W_ROM #(.FILENAME("conv11/CONV11_125.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U124 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(124+1)-1:16*124])); 
W_ROM #(.FILENAME("conv11/CONV11_126.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U125 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(125+1)-1:16*125])); 
W_ROM #(.FILENAME("conv11/CONV11_127.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U126 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(126+1)-1:16*126])); 
W_ROM #(.FILENAME("conv11/CONV11_128.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U127 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(127+1)-1:16*127])); 
W_ROM #(.FILENAME("conv11/CONV11_129.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U128 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(128+1)-1:16*128])); 
W_ROM #(.FILENAME("conv11/CONV11_130.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U129 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(129+1)-1:16*129])); 
W_ROM #(.FILENAME("conv11/CONV11_131.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U130 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(130+1)-1:16*130])); 
W_ROM #(.FILENAME("conv11/CONV11_132.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U131 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(131+1)-1:16*131])); 
W_ROM #(.FILENAME("conv11/CONV11_133.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U132 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(132+1)-1:16*132])); 
W_ROM #(.FILENAME("conv11/CONV11_134.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U133 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(133+1)-1:16*133])); 
W_ROM #(.FILENAME("conv11/CONV11_135.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U134 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(134+1)-1:16*134])); 
W_ROM #(.FILENAME("conv11/CONV11_136.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U135 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(135+1)-1:16*135])); 
W_ROM #(.FILENAME("conv11/CONV11_137.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U136 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(136+1)-1:16*136])); 
W_ROM #(.FILENAME("conv11/CONV11_138.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U137 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(137+1)-1:16*137])); 
W_ROM #(.FILENAME("conv11/CONV11_139.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U138 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(138+1)-1:16*138])); 
W_ROM #(.FILENAME("conv11/CONV11_140.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U139 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(139+1)-1:16*139])); 
W_ROM #(.FILENAME("conv11/CONV11_141.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U140 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(140+1)-1:16*140])); 
W_ROM #(.FILENAME("conv11/CONV11_142.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U141 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(141+1)-1:16*141])); 
W_ROM #(.FILENAME("conv11/CONV11_143.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U142 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(142+1)-1:16*142])); 
W_ROM #(.FILENAME("conv11/CONV11_144.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U143 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(143+1)-1:16*143])); 
W_ROM #(.FILENAME("conv11/CONV11_145.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U144 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(144+1)-1:16*144])); 
W_ROM #(.FILENAME("conv11/CONV11_146.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U145 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(145+1)-1:16*145])); 
W_ROM #(.FILENAME("conv11/CONV11_147.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U146 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(146+1)-1:16*146])); 
W_ROM #(.FILENAME("conv11/CONV11_148.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U147 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(147+1)-1:16*147])); 
W_ROM #(.FILENAME("conv11/CONV11_149.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U148 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(148+1)-1:16*148])); 
W_ROM #(.FILENAME("conv11/CONV11_150.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U149 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(149+1)-1:16*149])); 
W_ROM #(.FILENAME("conv11/CONV11_151.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U150 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(150+1)-1:16*150])); 
W_ROM #(.FILENAME("conv11/CONV11_152.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U151 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(151+1)-1:16*151])); 
W_ROM #(.FILENAME("conv11/CONV11_153.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U152 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(152+1)-1:16*152])); 
W_ROM #(.FILENAME("conv11/CONV11_154.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U153 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(153+1)-1:16*153])); 
W_ROM #(.FILENAME("conv11/CONV11_155.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U154 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(154+1)-1:16*154])); 
W_ROM #(.FILENAME("conv11/CONV11_156.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U155 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(155+1)-1:16*155])); 
W_ROM #(.FILENAME("conv11/CONV11_157.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U156 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(156+1)-1:16*156])); 
W_ROM #(.FILENAME("conv11/CONV11_158.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U157 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(157+1)-1:16*157])); 
W_ROM #(.FILENAME("conv11/CONV11_159.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U158 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(158+1)-1:16*158])); 
W_ROM #(.FILENAME("conv11/CONV11_160.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U159 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(159+1)-1:16*159])); 
W_ROM #(.FILENAME("conv11/CONV11_161.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U160 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(160+1)-1:16*160])); 
W_ROM #(.FILENAME("conv11/CONV11_162.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U161 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(161+1)-1:16*161])); 
W_ROM #(.FILENAME("conv11/CONV11_163.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U162 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(162+1)-1:16*162])); 
W_ROM #(.FILENAME("conv11/CONV11_164.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U163 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(163+1)-1:16*163])); 
W_ROM #(.FILENAME("conv11/CONV11_165.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U164 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(164+1)-1:16*164])); 
W_ROM #(.FILENAME("conv11/CONV11_166.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U165 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(165+1)-1:16*165])); 
W_ROM #(.FILENAME("conv11/CONV11_167.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U166 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(166+1)-1:16*166])); 
W_ROM #(.FILENAME("conv11/CONV11_168.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U167 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(167+1)-1:16*167])); 
W_ROM #(.FILENAME("conv11/CONV11_169.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U168 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(168+1)-1:16*168])); 
W_ROM #(.FILENAME("conv11/CONV11_170.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U169 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(169+1)-1:16*169])); 
W_ROM #(.FILENAME("conv11/CONV11_171.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U170 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(170+1)-1:16*170])); 
W_ROM #(.FILENAME("conv11/CONV11_172.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U171 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(171+1)-1:16*171])); 
W_ROM #(.FILENAME("conv11/CONV11_173.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U172 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(172+1)-1:16*172])); 
W_ROM #(.FILENAME("conv11/CONV11_174.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U173 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(173+1)-1:16*173])); 
W_ROM #(.FILENAME("conv11/CONV11_175.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U174 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(174+1)-1:16*174])); 
W_ROM #(.FILENAME("conv11/CONV11_176.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U175 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(175+1)-1:16*175])); 
W_ROM #(.FILENAME("conv11/CONV11_177.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U176 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(176+1)-1:16*176])); 
W_ROM #(.FILENAME("conv11/CONV11_178.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U177 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(177+1)-1:16*177])); 
W_ROM #(.FILENAME("conv11/CONV11_179.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U178 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(178+1)-1:16*178])); 
W_ROM #(.FILENAME("conv11/CONV11_180.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U179 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(179+1)-1:16*179])); 
W_ROM #(.FILENAME("conv11/CONV11_181.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U180 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(180+1)-1:16*180])); 
W_ROM #(.FILENAME("conv11/CONV11_182.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U181 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(181+1)-1:16*181])); 
W_ROM #(.FILENAME("conv11/CONV11_183.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U182 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(182+1)-1:16*182])); 
W_ROM #(.FILENAME("conv11/CONV11_184.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U183 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(183+1)-1:16*183])); 
W_ROM #(.FILENAME("conv11/CONV11_185.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U184 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(184+1)-1:16*184])); 
W_ROM #(.FILENAME("conv11/CONV11_186.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U185 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(185+1)-1:16*185])); 
W_ROM #(.FILENAME("conv11/CONV11_187.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U186 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(186+1)-1:16*186])); 
W_ROM #(.FILENAME("conv11/CONV11_188.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U187 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(187+1)-1:16*187])); 
W_ROM #(.FILENAME("conv11/CONV11_189.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U188 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(188+1)-1:16*188])); 
W_ROM #(.FILENAME("conv11/CONV11_190.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U189 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(189+1)-1:16*189])); 
W_ROM #(.FILENAME("conv11/CONV11_191.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U190 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(190+1)-1:16*190])); 
W_ROM #(.FILENAME("conv11/CONV11_192.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U191 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(191+1)-1:16*191])); 
W_ROM #(.FILENAME("conv11/CONV11_193.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U192 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(192+1)-1:16*192])); 
W_ROM #(.FILENAME("conv11/CONV11_194.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U193 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(193+1)-1:16*193])); 
W_ROM #(.FILENAME("conv11/CONV11_195.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U194 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(194+1)-1:16*194])); 
W_ROM #(.FILENAME("conv11/CONV11_196.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U195 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(195+1)-1:16*195])); 
W_ROM #(.FILENAME("conv11/CONV11_197.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U196 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(196+1)-1:16*196])); 
W_ROM #(.FILENAME("conv11/CONV11_198.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U197 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(197+1)-1:16*197])); 
W_ROM #(.FILENAME("conv11/CONV11_199.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U198 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(198+1)-1:16*198])); 
W_ROM #(.FILENAME("conv11/CONV11_200.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U199 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(199+1)-1:16*199])); 
W_ROM #(.FILENAME("conv11/CONV11_201.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U200 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(200+1)-1:16*200])); 
W_ROM #(.FILENAME("conv11/CONV11_202.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U201 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(201+1)-1:16*201])); 
W_ROM #(.FILENAME("conv11/CONV11_203.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U202 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(202+1)-1:16*202])); 
W_ROM #(.FILENAME("conv11/CONV11_204.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U203 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(203+1)-1:16*203])); 
W_ROM #(.FILENAME("conv11/CONV11_205.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U204 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(204+1)-1:16*204])); 
W_ROM #(.FILENAME("conv11/CONV11_206.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U205 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(205+1)-1:16*205])); 
W_ROM #(.FILENAME("conv11/CONV11_207.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U206 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(206+1)-1:16*206])); 
W_ROM #(.FILENAME("conv11/CONV11_208.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U207 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(207+1)-1:16*207])); 
W_ROM #(.FILENAME("conv11/CONV11_209.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U208 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(208+1)-1:16*208])); 
W_ROM #(.FILENAME("conv11/CONV11_210.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U209 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(209+1)-1:16*209])); 
W_ROM #(.FILENAME("conv11/CONV11_211.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U210 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(210+1)-1:16*210])); 
W_ROM #(.FILENAME("conv11/CONV11_212.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U211 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(211+1)-1:16*211])); 
W_ROM #(.FILENAME("conv11/CONV11_213.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U212 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(212+1)-1:16*212])); 
W_ROM #(.FILENAME("conv11/CONV11_214.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U213 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(213+1)-1:16*213])); 
W_ROM #(.FILENAME("conv11/CONV11_215.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U214 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(214+1)-1:16*214])); 
W_ROM #(.FILENAME("conv11/CONV11_216.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U215 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(215+1)-1:16*215])); 
W_ROM #(.FILENAME("conv11/CONV11_217.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U216 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(216+1)-1:16*216])); 
W_ROM #(.FILENAME("conv11/CONV11_218.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U217 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(217+1)-1:16*217])); 
W_ROM #(.FILENAME("conv11/CONV11_219.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U218 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(218+1)-1:16*218])); 
W_ROM #(.FILENAME("conv11/CONV11_220.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U219 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(219+1)-1:16*219])); 
W_ROM #(.FILENAME("conv11/CONV11_221.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U220 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(220+1)-1:16*220])); 
W_ROM #(.FILENAME("conv11/CONV11_222.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U221 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(221+1)-1:16*221])); 
W_ROM #(.FILENAME("conv11/CONV11_223.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U222 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(222+1)-1:16*222])); 
W_ROM #(.FILENAME("conv11/CONV11_224.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U223 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(223+1)-1:16*223])); 
W_ROM #(.FILENAME("conv11/CONV11_225.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U224 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(224+1)-1:16*224])); 
W_ROM #(.FILENAME("conv11/CONV11_226.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U225 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(225+1)-1:16*225])); 
W_ROM #(.FILENAME("conv11/CONV11_227.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U226 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(226+1)-1:16*226])); 
W_ROM #(.FILENAME("conv11/CONV11_228.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U227 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(227+1)-1:16*227])); 
W_ROM #(.FILENAME("conv11/CONV11_229.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U228 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(228+1)-1:16*228])); 
W_ROM #(.FILENAME("conv11/CONV11_230.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U229 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(229+1)-1:16*229])); 
W_ROM #(.FILENAME("conv11/CONV11_231.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U230 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(230+1)-1:16*230])); 
W_ROM #(.FILENAME("conv11/CONV11_232.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U231 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(231+1)-1:16*231])); 
W_ROM #(.FILENAME("conv11/CONV11_233.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U232 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(232+1)-1:16*232])); 
W_ROM #(.FILENAME("conv11/CONV11_234.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U233 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(233+1)-1:16*233])); 
W_ROM #(.FILENAME("conv11/CONV11_235.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U234 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(234+1)-1:16*234])); 
W_ROM #(.FILENAME("conv11/CONV11_236.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U235 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(235+1)-1:16*235])); 
W_ROM #(.FILENAME("conv11/CONV11_237.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U236 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(236+1)-1:16*236])); 
W_ROM #(.FILENAME("conv11/CONV11_238.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U237 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(237+1)-1:16*237])); 
W_ROM #(.FILENAME("conv11/CONV11_239.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U238 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(238+1)-1:16*238])); 
W_ROM #(.FILENAME("conv11/CONV11_240.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U239 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(239+1)-1:16*239])); 
W_ROM #(.FILENAME("conv11/CONV11_241.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U240 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(240+1)-1:16*240])); 
W_ROM #(.FILENAME("conv11/CONV11_242.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U241 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(241+1)-1:16*241])); 
W_ROM #(.FILENAME("conv11/CONV11_243.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U242 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(242+1)-1:16*242])); 
W_ROM #(.FILENAME("conv11/CONV11_244.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U243 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(243+1)-1:16*243])); 
W_ROM #(.FILENAME("conv11/CONV11_245.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U244 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(244+1)-1:16*244])); 
W_ROM #(.FILENAME("conv11/CONV11_246.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U245 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(245+1)-1:16*245])); 
W_ROM #(.FILENAME("conv11/CONV11_247.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U246 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(246+1)-1:16*246])); 
W_ROM #(.FILENAME("conv11/CONV11_248.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U247 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(247+1)-1:16*247])); 
W_ROM #(.FILENAME("conv11/CONV11_249.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U248 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(248+1)-1:16*248])); 
W_ROM #(.FILENAME("conv11/CONV11_250.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U249 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(249+1)-1:16*249])); 
W_ROM #(.FILENAME("conv11/CONV11_251.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U250 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(250+1)-1:16*250])); 
W_ROM #(.FILENAME("conv11/CONV11_252.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U251 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(251+1)-1:16*251])); 
W_ROM #(.FILENAME("conv11/CONV11_253.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U252 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(252+1)-1:16*252])); 
W_ROM #(.FILENAME("conv11/CONV11_254.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U253 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(253+1)-1:16*253])); 
W_ROM #(.FILENAME("conv11/CONV11_255.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U254 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(254+1)-1:16*254])); 
W_ROM #(.FILENAME("conv11/CONV11_256.txt"),.weight_addr_WIDTH(3),.NO_ROWS(7)) U255 (.weight_addr(weight_addr_conv11),.clk(clk),.weight_out(weight_out_conv11[16*(255+1)-1:16*255])); 


endmodule

