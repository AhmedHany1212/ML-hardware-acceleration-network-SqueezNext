module BIAS_L2 #(parameter N=48)(out,Z,U);
wire [N*18-1:0] q;
input Z,U;
output reg [N/3*18-1:0] out;

always @(*)
begin
	case({U,Z})
		2'b10: out=q[18*16-1:18*0];
		2'b11: out=q[18*32-1:18*16];
		2'b00: out=q[18*48-1:18*32];
		default:out=0;
	endcase
end

BIAS #(.value(18'b000001111110100000)) U0 (.q(q[18*(0+1)-1:18*0])); 
BIAS #(.value(18'b111101101010011000)) U1 (.q(q[18*(1+1)-1:18*1])); 
BIAS #(.value(18'b000001100010011000)) U2 (.q(q[18*(2+1)-1:18*2])); 
BIAS #(.value(18'b001001101101100000)) U3 (.q(q[18*(3+1)-1:18*3])); 
BIAS #(.value(18'b001000101111110000)) U4 (.q(q[18*(4+1)-1:18*4])); 
BIAS #(.value(18'b000001011011000000)) U5 (.q(q[18*(5+1)-1:18*5])); 
BIAS #(.value(18'b111111101100001000)) U6 (.q(q[18*(6+1)-1:18*6])); 
BIAS #(.value(18'b111111000010110100)) U7 (.q(q[18*(7+1)-1:18*7])); 
BIAS #(.value(18'b000001001000101100)) U8 (.q(q[18*(8+1)-1:18*8])); 
BIAS #(.value(18'b000000110110011000)) U9 (.q(q[18*(9+1)-1:18*9])); 
BIAS #(.value(18'b000010110111100000)) U10 (.q(q[18*(10+1)-1:18*10])); 
BIAS #(.value(18'b111111110001000000)) U11 (.q(q[18*(11+1)-1:18*11])); 
BIAS #(.value(18'b000100010010011000)) U12 (.q(q[18*(12+1)-1:18*12])); 
BIAS #(.value(18'b000001100100010100)) U13 (.q(q[18*(13+1)-1:18*13])); 
BIAS #(.value(18'b111101000010011100)) U14 (.q(q[18*(14+1)-1:18*14])); 
BIAS #(.value(18'b111111111100100000)) U15 (.q(q[18*(15+1)-1:18*15]));
 
BIAS #(.value(18'b000100100000101100)) U16 (.q(q[18*(16+1)-1:18*16])); 
BIAS #(.value(18'b111111011001100000)) U17 (.q(q[18*(17+1)-1:18*17])); 
BIAS #(.value(18'b000010110110000100)) U18 (.q(q[18*(18+1)-1:18*18])); 
BIAS #(.value(18'b000010000111111100)) U19 (.q(q[18*(19+1)-1:18*19])); 
BIAS #(.value(18'b111111111110000000)) U20 (.q(q[18*(20+1)-1:18*20])); 
BIAS #(.value(18'b111111111100010000)) U21 (.q(q[18*(21+1)-1:18*21])); 
BIAS #(.value(18'b000101011001101000)) U22 (.q(q[18*(22+1)-1:18*22])); 
BIAS #(.value(18'b000010110001101000)) U23 (.q(q[18*(23+1)-1:18*23])); 
BIAS #(.value(18'b111011110011001000)) U24 (.q(q[18*(24+1)-1:18*24])); 
BIAS #(.value(18'b000110111010110100)) U25 (.q(q[18*(25+1)-1:18*25])); 
BIAS #(.value(18'b000101000001110000)) U26 (.q(q[18*(26+1)-1:18*26])); 
BIAS #(.value(18'b111110010101001100)) U27 (.q(q[18*(27+1)-1:18*27])); 
BIAS #(.value(18'b111111011110000100)) U28 (.q(q[18*(28+1)-1:18*28])); 
BIAS #(.value(18'b111101101100010000)) U29 (.q(q[18*(29+1)-1:18*29])); 
BIAS #(.value(18'b000001101010111100)) U30 (.q(q[18*(30+1)-1:18*30])); 
BIAS #(.value(18'b111111001101110000)) U31 (.q(q[18*(31+1)-1:18*31])); 

BIAS #(.value(18'b000000001001111100)) U32 (.q(q[18*(32+1)-1:18*32])); 
BIAS #(.value(18'b111110010100111000)) U33 (.q(q[18*(33+1)-1:18*33])); 
BIAS #(.value(18'b001011011000011100)) U34 (.q(q[18*(34+1)-1:18*34])); 
BIAS #(.value(18'b000110101111011000)) U35 (.q(q[18*(35+1)-1:18*35])); 
BIAS #(.value(18'b110110111010101000)) U36 (.q(q[18*(36+1)-1:18*36])); 
BIAS #(.value(18'b000101011000011000)) U37 (.q(q[18*(37+1)-1:18*37])); 
BIAS #(.value(18'b000010101100110000)) U38 (.q(q[18*(38+1)-1:18*38])); 
BIAS #(.value(18'b111101000111111100)) U39 (.q(q[18*(39+1)-1:18*39])); 
BIAS #(.value(18'b111011110100100000)) U40 (.q(q[18*(40+1)-1:18*40])); 
BIAS #(.value(18'b111111001001100000)) U41 (.q(q[18*(41+1)-1:18*41])); 
BIAS #(.value(18'b000110010110100100)) U42 (.q(q[18*(42+1)-1:18*42])); 
BIAS #(.value(18'b001000010010100000)) U43 (.q(q[18*(43+1)-1:18*43])); 
BIAS #(.value(18'b111111101111101100)) U44 (.q(q[18*(44+1)-1:18*44])); 
BIAS #(.value(18'b000001111100100100)) U45 (.q(q[18*(45+1)-1:18*45])); 
BIAS #(.value(18'b000001001010000000)) U46 (.q(q[18*(46+1)-1:18*46])); 
BIAS #(.value(18'b111111100111010000)) U47 (.q(q[18*(47+1)-1:18*47])); 

endmodule